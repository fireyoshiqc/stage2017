use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

library work;
use work.util.all;

entity system is
port(
    start : in std_logic;
    test_out : out std_logic_vector(8 - 1 downto 0);
    sel : in unsigned(8 - 1 downto 0)
);
end system;

architecture system of system is

component fc_layer is
generic(
    input_width : integer;
    output_width : integer;
    simd_width : integer;
    input_spec : fixed_spec;
    weight_spec : fixed_spec;
    op_arg_spec : fixed_spec;
    output_spec : fixed_spec;
    n_weights : integer;
    weights_filename : string;
    weight_values : reals
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    in_a : in std_logic_vector;
    out_a : out std_logic_vector;
    out_offset : out unsigned;
    op_argument : out sfixed;
    op_result : in sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component interlayer is
generic(
    width : integer;
    word_size : integer
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    ack : out std_logic;
    previous_a : in std_logic_vector;
    next_a : out std_logic_vector
);
end component;

component bias_op is
generic(
    input_spec : fixed_spec;
    bias_spec : fixed_spec;
    biases : reals
);
port(
    input : in sfixed;
    offset : in unsigned;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component sigmoid_op is
generic(
    input_spec : fixed_spec;
    output_spec : fixed_spec;
    step_precision : integer;
    bit_precision : integer
);
port(
    clk : in std_logic;
    input : in sfixed;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;




signal ready_s1 : std_logic;
signal done_s2 : std_logic;
signal start_s3 : std_logic;
signal ack_s4 : std_logic;
signal in_a_s5 : std_logic_vector(7055 downto 0);
signal out_a_s6 : std_logic_vector(399 downto 0);
signal out_offset_s7 : unsigned(5 downto 0);
signal op_argument_s8 : sfixed(13 downto -14);
signal op_result_s9 : sfixed(1 downto -8);
signal op_send_s10 : std_logic;
signal op_receive_s11 : std_logic;



signal ready_s71 : std_logic;
signal done_s72 : std_logic;
signal start_s73 : std_logic;
signal ack_s74 : std_logic;
signal previous_a_s75 : std_logic_vector(7055 downto 0);
signal next_a_s76 : std_logic_vector(7055 downto 0);

signal input_s13 : sfixed(13 downto -14);
signal offset_s14 : unsigned(5 downto 0);
signal output_s15 : sfixed(14 downto -14);
signal op_send_s16 : std_logic;
signal op_receive_s17 : std_logic;


signal input_s19 : sfixed(14 downto -14);
signal output_s20 : sfixed(1 downto -8);
signal op_send_s21 : std_logic;
signal op_receive_s22 : std_logic;



signal ready_s24 : std_logic;
signal done_s25 : std_logic;
signal start_s26 : std_logic;
signal ack_s27 : std_logic;
signal in_a_s28 : std_logic_vector(399 downto 0);
signal out_a_s29 : std_logic_vector(399 downto 0);
signal out_offset_s30 : unsigned(5 downto 0);
signal op_argument_s31 : sfixed(12 downto -13);
signal op_result_s32 : sfixed(1 downto -8);
signal op_send_s33 : std_logic;
signal op_receive_s34 : std_logic;



signal ready_s95 : std_logic;
signal done_s96 : std_logic;
signal start_s97 : std_logic;
signal ack_s98 : std_logic;
signal previous_a_s99 : std_logic_vector(399 downto 0);
signal next_a_s100 : std_logic_vector(399 downto 0);

signal input_s36 : sfixed(12 downto -13);
signal offset_s37 : unsigned(5 downto 0);
signal output_s38 : sfixed(13 downto -13);
signal op_send_s39 : std_logic;
signal op_receive_s40 : std_logic;


signal input_s42 : sfixed(13 downto -13);
signal output_s43 : sfixed(1 downto -8);
signal op_send_s44 : std_logic;
signal op_receive_s45 : std_logic;



signal ready_s47 : std_logic;
signal done_s48 : std_logic;
signal start_s49 : std_logic;
signal ack_s50 : std_logic;
signal in_a_s51 : std_logic_vector(399 downto 0);
signal out_a_s52 : std_logic_vector(99 downto 0);
signal out_offset_s53 : unsigned(3 downto 0);
signal op_argument_s54 : sfixed(13 downto -12);
signal op_result_s55 : sfixed(1 downto -8);
signal op_send_s56 : std_logic;
signal op_receive_s57 : std_logic;



signal ready_s103 : std_logic;
signal done_s104 : std_logic;
signal start_s105 : std_logic;
signal ack_s106 : std_logic;
signal previous_a_s107 : std_logic_vector(399 downto 0);
signal next_a_s108 : std_logic_vector(399 downto 0);

signal input_s59 : sfixed(13 downto -12);
signal offset_s60 : unsigned(3 downto 0);
signal output_s61 : sfixed(14 downto -12);
signal op_send_s62 : std_logic;
signal op_receive_s63 : std_logic;


signal input_s65 : sfixed(14 downto -12);
signal output_s66 : sfixed(1 downto -8);
signal op_send_s67 : std_logic;
signal op_receive_s68 : std_logic;


component ps is
port(
    clk, rst : out std_logic
);
end component;

signal clk, rst_sink : std_logic;
constant rst : std_logic := '0';

function to_vec(r : reals) return std_logic_vector is
    constant input_spec : fixed_spec := fixed_spec(fixed_spec'(int => 1, frac => 8));
    variable ret : std_logic_vector(784 * size(input_spec) - 1 downto 0);
begin
    for i in r'range loop
        ret((1 + i) * size(input_spec) - 1 downto i * size(input_spec)) :=
            std_logic_vector(to_sfixed(r(i), mk(input_spec)));
    end loop;
    return ret;
end to_vec;

begin

fc_layer_u0 : fc_layer generic map(
    input_width => 784,
    output_width => 40,
    simd_width => 14,
    input_spec => fixed_spec(fixed_spec'(int => 1, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 2, frac => 6)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 14, frac => 14)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    n_weights => 31360,
    weights_filename => "whatever",
    weight_values => reals(reals'( 0.0000408, 0.0001156, -0.0007705, -0.0003351, -0.0000950, -0.0000820, 0.0004032, 0.0004182, 0.0003001, -0.0001907, 0.0000297, 0.0001292, 0.0016181, 0.0033509, -0.0004116, 0.0003559, -0.0004802, 0.0006479, 0.0000861, 0.0001580, -0.0002336, -0.0007931, 0.0001428, 0.0002428, 0.0001890, 0.0001554, 0.0000769, -0.0002156, -0.0003911, 0.0005581, -0.0002465, 0.0002428, -0.0002677, 0.0001292, 0.0038330, 0.0061119, 0.0063058, 0.0006660, 0.0018109, 0.0006858, 0.0013706, -0.0008381, -0.0072303, -0.0185001, -0.0347154, -0.0061202, 0.0011924, 0.0005082, 0.0053583, 0.0091062, 0.0035945, 0.0034690, -0.0000003, -0.0001222, -0.0000568, 0.0004877, -0.0001252, 0.0003127, -0.0004140, -0.0001421, -0.0000033, 0.0006630, 0.0109417, 0.0252189, 0.0151279, 0.0068338, 0.0396617, 0.0650002, 0.0643596, 0.0811151, 0.0860193, -0.0110326, -0.0857354, -0.0706970, -0.0742991, -0.0005925, 0.0023063, 0.0138023, 0.0146258, 0.0043074, 0.0012573, -0.0001469, 0.0000623, 0.0000403, -0.0004547, -0.0000152, -0.0005816, -0.0001612, -0.0031084, 0.0046655, 0.0184095, 0.0547722, 0.0458653, 0.0764468, 0.0815437, 0.1466200, 0.0937492, 0.0375963, 0.0035690, -0.1021800, -0.2487210, -0.3082000, -0.2899820, -0.0337810, 0.0001316, 0.0216308, 0.0618042, 0.0580215, 0.0566176, 0.0078293, 0.0029489, 0.0002086, 0.0003119, 0.0001715, -0.0005010, -0.0004678, 0.0152223, 0.0533587, 0.0362833, 0.0299187, 0.0700633, 0.0895389, 0.1649460, 0.1331820, 0.1819780, 0.0565010, -0.1609890, -0.4032590, -0.4190330, -0.3572230, -0.1928310, 0.0605936, 0.0882286, 0.0867366, 0.1055950, 0.0875757, -0.0268386, -0.0430774, -0.0172364, 0.0036921, 0.0001532, 0.0001673, -0.0000059, -0.0072398, 0.0208059, 0.1688750, 0.1909760, 0.0865629, 0.1039180, 0.2798850, 0.3238080, 0.1378940, 0.2829040, -0.2263370, -0.6018320, -0.8534070, -0.5163420, -0.0100411, 0.1574760, 0.2480940, 0.0461678, 0.0378534, 0.0724771, 0.1342370, 0.0580798, -0.0394766, 0.0024487, 0.0076129, 0.0000928, 0.0003728, -0.0064206, -0.0605344, -0.0266544, 0.1227010, 0.1451860, 0.1449620, 0.2019420, 0.2780500, 0.1807230, 0.2340500, 0.1263620, -0.1964740, -0.9113080, -1.1540300, -0.4700730, 0.0665744, 0.1417590, 0.2358060, 0.1873120, -0.0416665, 0.0090010, 0.1549920, 0.0240485, -0.0267736, 0.0006723, 0.0077243, -0.0000285, 0.0023462, -0.0025640, -0.0657071, -0.0152877, 0.0693240, 0.0630817, 0.0741730, 0.0615562, 0.2631320, 0.3346370, 0.2321780, -0.0041563, -0.3724530, -0.8663880, -0.8247520, -0.2379330, 0.0877544, 0.1769310, 0.2037680, 0.1364920, 0.0265569, 0.0691599, 0.0900181, -0.1163740, -0.0665033, 0.0174623, 0.0040099, 0.0009015, 0.0038694, 0.0061569, -0.0065498, 0.0100425, 0.0665915, 0.0086675, 0.1650280, 0.1150910, 0.2559440, 0.2103880, 0.3606190, 0.3568610, -0.2033450, -0.8553220, -0.5303120, 0.0843481, 0.2036230, 0.1661590, 0.1818670, -0.0499374, -0.0155624, -0.0014863, -0.0768179, -0.1490330, -0.0253135, -0.0357896, -0.0058015, -0.0002553, 0.0029923, 0.0110067, 0.0237443, 0.0846660, 0.0344682, -0.0391484, 0.0321596, 0.2034950, 0.0690879, 0.0916413, 0.3515740, 0.4030360, -0.3933870, -0.8713900, -0.0857388, 0.3325590, 0.2552340, 0.1656670, 0.1179140, 0.0361244, 0.0444135, 0.0276070, -0.0936895, -0.0007871, -0.0660689, -0.0471792, 0.0069456, 0.0001135, 0.0033795, 0.0222199, 0.0046883, 0.1319100, 0.0727055, -0.2025440, -0.0965611, 0.1306940, 0.0372889, 0.0024322, 0.3224870, 0.1386070, -0.7207660, -0.6768400, -0.0494575, 0.2243560, 0.2467750, 0.0564180, 0.1677640, -0.0048336, 0.1933900, 0.0008101, -0.0728858, 0.0831703, 0.0314235, -0.0194856, -0.0025027, 0.0003479, 0.0041175, 0.0050364, -0.0131561, 0.0649843, 0.0597026, -0.1620470, -0.2529410, -0.1225150, -0.2856400, -0.1759120, -0.0267279, -0.1076350, -0.4435970, -0.0710733, -0.0131802, 0.1068500, 0.0843650, 0.1885230, -0.0146504, -0.0342709, 0.1375340, -0.0521685, -0.0173079, 0.0171801, 0.0077618, -0.0231124, -0.0034051, 0.0001255, 0.0022242, 0.0204442, -0.0053252, 0.0119030, -0.0699116, -0.0808024, -0.0198391, -0.0490748, -0.3275890, -0.0885521, -0.0497274, -0.2151700, -0.2163290, -0.0213713, 0.1578520, 0.2068590, 0.1116020, -0.0059451, -0.0894573, 0.0617414, 0.1435130, 0.0796905, 0.0125305, 0.1085390, 0.0247227, -0.0277629, -0.0024571, -0.0003229, 0.0012920, 0.0103546, -0.0106631, -0.0164188, -0.0568550, 0.0814357, 0.0269486, -0.1084900, -0.1312440, -0.0582799, -0.1737650, -0.1614230, -0.1084430, -0.1222190, 0.0547736, 0.0218422, 0.1035710, 0.0505919, 0.0172878, 0.1239620, 0.0842178, 0.0065643, 0.1280380, 0.1073900, 0.0033204, -0.0505904, -0.0089756, -0.0004512, 0.0007733, 0.0088420, 0.0046793, -0.0745362, 0.0867803, -0.0288933, -0.0898602, -0.1502590, -0.0455147, -0.0503216, -0.0765177, -0.1034450, 0.0344278, 0.0892354, 0.0600338, 0.1526920, 0.1840780, -0.0668432, 0.2106850, 0.0314651, 0.0917470, 0.1516250, 0.1599450, 0.0597286, -0.0562202, -0.0456400, -0.0007958, -0.0009939, -0.0001021, -0.0059756, 0.0059784, -0.1118230, -0.1156010, -0.0295223, -0.0486842, -0.0676776, -0.0418525, -0.0477763, -0.1402360, -0.0615344, 0.1774690, 0.0716666, 0.0875325, -0.0136577, 0.0199230, -0.1230670, -0.0388063, -0.0305183, 0.0591164, 0.1687850, 0.0557864, -0.0905482, -0.0750084, -0.0004287, -0.0021150, 0.0001570, -0.0004730, -0.0298011, -0.0402610, -0.1746850, -0.1948710, -0.0762271, -0.1859970, 0.0100104, 0.0141201, -0.0622938, -0.0950794, 0.1562120, 0.0405879, 0.1078830, 0.1261290, 0.1046360, -0.0174896, 0.0889589, 0.0474537, -0.0515373, 0.0813138, -0.0744943, -0.0717250, -0.0936186, -0.0444926, -0.0427723, -0.0035386, -0.0002195, 0.0006087, -0.0325336, -0.0951248, -0.1684800, -0.1524870, -0.0364741, -0.1845130, -0.0957929, 0.0254724, 0.0736886, 0.1413140, 0.0382526, -0.1458960, 0.1215090, 0.0214734, 0.1577360, 0.0706191, 0.1519460, -0.0324796, -0.2222560, -0.0485154, 0.0112820, 0.0962036, 0.0518066, 0.0549371, -0.0092330, -0.0106889, -0.0007506, -0.0004864, -0.0048412, -0.0878337, -0.2129410, -0.2382620, -0.2094190, 0.0235527, 0.0458034, 0.0668059, -0.0421649, 0.1480100, -0.0571565, -0.0349147, 0.0603500, 0.1080350, -0.0681785, 0.1111850, -0.0295117, -0.1629920, -0.2659610, -0.0957737, 0.0463551, 0.1180560, 0.0327841, 0.0305466, -0.0030399, -0.0026610, 0.0002386, -0.0002915, -0.0020334, -0.0273103, -0.2076640, -0.2611830, -0.1460090, -0.0140140, -0.0036005, -0.0221827, 0.0293505, 0.0965633, -0.1817490, -0.0730674, 0.0356824, 0.1392200, 0.0053140, -0.0389051, -0.2184490, -0.1581750, -0.0966867, -0.0971920, -0.0688112, 0.0289225, -0.0425716, -0.0111752, -0.0014794, -0.0002943, 0.0002747, -0.0002694, -0.0034933, -0.0403083, -0.1096950, -0.3176500, -0.0881138, 0.0417062, -0.0558304, -0.1053110, -0.1244970, -0.0864638, -0.0600173, -0.0991870, 0.0108096, 0.0973347, 0.1477070, 0.0050927, 0.0448658, -0.0700960, -0.0826448, -0.0806831, -0.0461665, 0.0122476, -0.0856628, -0.0543442, -0.0008070, -0.0004491, 0.0003790, 0.0001805, -0.0047105, -0.0223951, -0.0364490, 0.0540679, 0.1183840, 0.1417220, 0.2007610, -0.0518821, -0.0669496, -0.0036837, -0.0570206, 0.0368226, -0.0216283, -0.0309799, 0.0519017, 0.0853929, -0.0738333, -0.1757540, 0.0094682, -0.0165018, -0.0800523, 0.0231095, 0.0036233, -0.0263544, 0.0006321, 0.0006996, -0.0002790, 0.0006154, 0.0005682, -0.0258020, 0.0293326, 0.1470070, 0.1084000, -0.0077538, 0.1534960, 0.1394860, -0.0098732, -0.0139355, -0.1278760, 0.0582982, -0.1863740, -0.0114817, 0.0433498, -0.0455971, -0.1169080, -0.0058821, -0.0736090, -0.0709483, -0.0807464, -0.1099060, -0.0353974, -0.0025672, 0.0083444, -0.0002610, -0.0000219, 0.0004906, -0.0063589, -0.0435964, -0.0490502, -0.0356928, -0.0509430, 0.0111657, 0.0109166, 0.0396625, 0.1332030, -0.0957493, -0.0085857, 0.0457823, -0.1557700, -0.1246830, -0.0348519, -0.0693903, -0.0997581, -0.0158861, -0.1263150, -0.1260530, -0.1406870, -0.1419620, -0.0784485, 0.0178957, 0.0088947, 0.0005972, 0.0000757, -0.0000196, -0.0079887, -0.0129567, -0.0468040, -0.0374206, -0.1315180, -0.1116230, -0.0516431, -0.0143117, -0.0163546, 0.0047835, 0.0603702, 0.3281290, 0.1504540, 0.0503262, 0.0671761, 0.0084153, 0.0184817, -0.1537120, -0.2056200, -0.1279210, -0.1163730, -0.0822051, -0.0366765, -0.0015442, 0.0000140, 0.0002774, 0.0002554, -0.0000816, -0.0019452, 0.0030543, -0.0265426, -0.0331130, -0.0933214, -0.0953786, 0.0157823, -0.0912639, -0.0913371, 0.0716800, 0.0861137, 0.0629052, 0.0565487, -0.0249400, 0.0419544, -0.0404942, -0.0745949, -0.2468560, -0.1708230, -0.1106010, -0.0481797, 0.0135830, -0.0036545, 0.0000869, 0.0005060, 0.0001490, 0.0001019, -0.0003215, 0.0004246, -0.0002209, -0.0016589, -0.0462476, -0.0743337, -0.0679151, -0.0720385, -0.0810903, -0.1314830, -0.1473480, -0.1723090, -0.1391910, -0.1182880, 0.0058996, 0.0481091, -0.0290945, -0.0273430, -0.0258332, -0.0547328, -0.0708932, -0.0268237, -0.0098079, -0.0017526, 0.0001125, 0.0002152, -0.0003248, -0.0002191, -0.0003299, -0.0001119, 0.0002347, 0.0005113, 0.0012863, 0.0000768, -0.0104565, -0.0076258, 0.0067648, 0.0143351, 0.0033226, 0.0089187, 0.0286165, -0.0142253, -0.0110749, -0.0029500, -0.0035345, -0.0403840, -0.0145956, -0.0054587, -0.0053104, -0.0132141, -0.0001621, -0.0002462, -0.0000518, 0.0003005, 0.0005547, 0.0005017, 0.0003417, 0.0005156, -0.0005799, -0.0003289, 0.0003080, 0.0002153, -0.0002026, -0.0005443, -0.0000155, -0.0002491, -0.0000362, 0.0008848, 0.0004049, -0.0002092, -0.0000238, -0.0001995, -0.0004874, -0.0003552, -0.0003460, 0.0000113, 0.0005768, -0.0005318, -0.0000948, -0.0003511, 0.0000383, 0.0001099, 0.0000532, -0.0004529, -0.0001624, 0.0004796, 0.0000320, 0.0001740, 0.0000467, 0.0003068, 0.0000069, -0.0000238, -0.0001619, -0.0016537, -0.0063152, -0.0002852, 0.0011523, 0.0087804, 0.0448993, 0.0334157, 0.0160667, 0.0046870, 0.0117603, 0.0187377, 0.0156275, 0.0012687, 0.0000278, 0.0002506, 0.0001123, -0.0000300, 0.0002314, -0.0000043, -0.0000965, -0.0000811, 0.0009823, 0.0014335, 0.0001440, 0.0002692, 0.0001640, -0.0005229, -0.0031788, -0.0215140, -0.0332750, 0.0096054, -0.0249847, -0.0396970, 0.0039847, 0.0026207, -0.0073925, 0.0748362, 0.0489993, 0.0174990, -0.0011929, -0.0007676, 0.0036706, 0.0017560, 0.0004104, 0.0001484, -0.0003306, -0.0003661, 0.0007411, 0.0002006, 0.0038785, 0.0037628, -0.0005562, -0.0012528, -0.0011835, -0.0231292, -0.0287376, -0.0309792, -0.1068680, -0.0504197, -0.0782426, -0.0509338, 0.0130941, -0.0150066, 0.0585860, 0.1713180, 0.0602553, 0.0579530, -0.0215167, 0.0056434, 0.0048402, -0.0022889, 0.0272559, 0.0081389, -0.0002473, -0.0003850, 0.0007205, 0.0000037, 0.0001276, 0.0031170, 0.0036788, -0.0030590, -0.0311929, -0.0992892, -0.2277340, -0.2860040, -0.2107680, -0.2315490, -0.1363720, -0.0187810, 0.0379730, 0.0573720, -0.0760982, -0.0856629, 0.0588856, -0.0055431, 0.0219984, 0.0934437, 0.1132700, 0.0694466, 0.0408566, 0.0122362, 0.0012939, 0.0001742, 0.0001716, -0.0002143, 0.0028698, 0.0545935, 0.1133830, 0.0686728, 0.0085953, -0.0619862, -0.0381337, -0.0898982, -0.1776430, -0.2120530, 0.1015030, 0.0716205, -0.0427944, -0.1482060, -0.0301596, -0.1442570, -0.0753183, 0.0576598, -0.1258830, -0.0494794, 0.0028584, 0.0442150, 0.0284218, 0.0164900, -0.0010766, 0.0005644, -0.0000432, 0.0012568, 0.0192511, 0.0769439, 0.0617554, 0.0281946, -0.0274883, -0.0700405, -0.1857980, -0.0524282, -0.2036400, -0.1536910, 0.0192214, -0.0518016, 0.0393519, 0.0554600, 0.0929111, 0.1703130, 0.1057390, 0.2013160, 0.0187339, -0.0493770, -0.0733107, -0.0047502, 0.0350211, 0.0256373, -0.0006927, 0.0000951, -0.0008204, -0.0033538, 0.0392777, 0.0419978, -0.0259616, -0.0637981, -0.0867003, -0.2724920, -0.2444630, -0.1365910, -0.2290580, 0.1503310, -0.1908370, -0.0905033, 0.0854404, 0.2828320, 0.3552940, 0.1678900, 0.1827300, 0.1946530, 0.0358451, 0.0039315, 0.0719386, -0.0745950, 0.0011671, 0.0274306, 0.0015518, 0.0015090, -0.0015635, 0.0053774, 0.0444339, 0.0022789, 0.0080412, -0.0233302, -0.0839905, -0.1994180, -0.2102080, -0.2116520, -0.2379260, -0.0850184, -0.1333760, -0.1326680, 0.1183300, 0.4423790, 0.3640090, 0.1984620, -0.0199276, 0.0297248, 0.1205210, 0.1107310, -0.0267557, 0.0074573, -0.0006575, 0.0416149, 0.0058837, 0.0003265, 0.0033472, 0.0059062, 0.0154411, 0.0337434, 0.0340231, 0.0185949, -0.1432860, -0.1053910, -0.1030680, -0.1395610, -0.1085750, 0.1165330, -0.0685289, -0.1559360, -0.0083870, 0.1482710, 0.2338760, 0.0065076, 0.0882311, 0.1040850, 0.0750237, 0.2003660, 0.0309338, 0.1164320, 0.1541700, 0.0460717, 0.0180476, 0.0004022, 0.0007973, 0.0215506, -0.0070523, 0.0717181, -0.0115780, -0.1115840, -0.1469990, -0.0883728, -0.1438380, -0.0145118, 0.1117780, -0.0372669, -0.0053898, 0.0186662, -0.0151516, 0.2069600, -0.0097955, 0.1197930, 0.1829240, 0.2469160, 0.0280067, 0.2262600, 0.1849240, 0.1631070, 0.0940779, 0.0083726, 0.0032828, 0.0003528, 0.0032978, 0.0165420, 0.0007371, 0.0124750, -0.0531904, -0.1010700, 0.0492094, -0.0462765, -0.1243920, -0.0025783, -0.0172913, -0.1748070, 0.1309550, 0.2766660, 0.0265647, -0.0764470, 0.1882590, 0.2928750, 0.2552080, 0.3012690, 0.2375540, 0.1964010, 0.1900410, 0.1676910, 0.0166030, 0.0125277, 0.0015314, -0.0000888, 0.0003142, 0.0043521, 0.0017417, -0.0153591, -0.0454617, -0.0972373, -0.0916195, -0.1882540, 0.0140081, -0.0175148, -0.0716265, -0.2756710, -0.1465130, 0.2734660, 0.1532760, -0.1043600, 0.0179967, 0.1595770, 0.1491590, 0.0009187, -0.1258110, 0.0901275, 0.1842600, -0.0163937, -0.0266343, 0.0095632, 0.0036485, 0.0005293, -0.0001503, 0.0013842, 0.0046433, 0.0632242, -0.0517690, -0.1577180, -0.2196990, -0.1031490, -0.0569945, -0.1367410, -0.1422990, -0.1751280, -0.0653755, 0.1310640, 0.0833074, -0.0470368, -0.1310010, -0.1609580, -0.0904492, -0.1136490, -0.0919171, -0.0271961, -0.0774207, -0.0835079, -0.0350975, -0.0225090, -0.0030900, 0.0002240, 0.0010612, 0.0001466, 0.0064878, 0.0086235, -0.0368759, -0.0722270, -0.1748210, -0.0543359, -0.1652430, -0.0341593, -0.2289210, -0.2613350, -0.0576424, 0.0348660, 0.0440127, -0.2284620, -0.2461160, -0.2726630, -0.1127890, 0.0460345, -0.0307470, -0.2324520, -0.1705740, -0.0741004, -0.0577297, -0.0114036, -0.0001884, -0.0002182, 0.0004218, -0.0045453, -0.0505959, 0.0366973, 0.0346020, 0.1157000, 0.1075580, -0.1336870, -0.2767180, -0.0373944, -0.1780870, -0.1079740, -0.0752217, -0.0740654, 0.1312290, -0.0390551, -0.1316060, -0.1701290, -0.1037890, -0.1026570, -0.2761280, -0.2033650, -0.0871825, -0.0811728, -0.0581286, -0.0198657, -0.0039295, 0.0003116, 0.0007488, -0.0160391, -0.0824786, 0.0661951, 0.1217300, 0.1549450, -0.0269492, -0.0684621, -0.0918685, 0.0919643, -0.2209800, -0.1025780, -0.1168660, -0.2745330, -0.0911390, 0.1747660, -0.1485390, -0.1510300, -0.1332750, -0.2422400, -0.4066150, -0.2736420, -0.2472390, -0.0983226, -0.0653812, -0.0202670, -0.0019405, 0.0007615, 0.0000556, -0.0411603, -0.0790447, -0.0611755, 0.0371314, -0.0218837, 0.0741209, -0.0946739, -0.0266463, -0.0687393, -0.0676540, -0.0439938, -0.1281180, -0.0152750, 0.0401833, 0.3409900, 0.1735750, -0.0077868, -0.1368260, -0.3555340, -0.4474650, -0.2647700, -0.0837455, -0.0323890, -0.0093414, -0.0003000, 0.0034934, 0.0020195, 0.0001020, -0.0113652, -0.1255090, -0.0942642, 0.0438403, -0.1168460, -0.0631393, -0.0984136, -0.0157351, 0.0042044, 0.1948170, 0.0701502, 0.0271352, 0.0024219, 0.2316930, 0.4222540, 0.3713020, 0.0465020, -0.4545460, -0.5087490, -0.4268030, -0.2510450, -0.1740120, -0.0937996, 0.0003356, 0.0018239, -0.0031458, -0.0000154, 0.0130576, 0.0101637, -0.0705998, -0.1049480, 0.0056424, 0.0551895, -0.0408438, -0.0521595, -0.0393593, -0.0083495, -0.0510184, 0.1000240, 0.0028206, 0.1309820, 0.0648546, 0.2699960, 0.3166940, -0.0836456, -0.6341840, -0.4372990, -0.2974070, -0.1514620, -0.1006770, 0.0097033, 0.0319331, -0.0062322, -0.0007719, 0.0000388, 0.0047803, 0.0014365, -0.0493511, -0.1017720, -0.0378380, 0.0623866, -0.1078000, -0.0128991, 0.0145021, 0.1347020, 0.0556604, 0.0574085, 0.1091950, -0.0369700, 0.0784687, 0.0277079, 0.2193850, -0.5216880, -0.8209180, -0.5295420, -0.2371090, -0.0593632, -0.0714507, 0.0126953, 0.0151494, -0.0036670, -0.0000233, 0.0003118, -0.0005654, -0.0074893, -0.0514320, -0.1726690, -0.1969270, -0.0189953, 0.0328367, 0.0380959, 0.0156400, 0.0724502, -0.0442976, -0.0389969, -0.1818740, -0.0147908, 0.0000416, -0.1401650, -0.2048130, -0.6952940, -0.6081020, -0.3082100, -0.1093220, -0.0586622, -0.0377498, -0.0161735, -0.0003245, 0.0059131, 0.0003303, 0.0002252, 0.0000185, -0.0071507, -0.0424889, -0.1251670, -0.1659400, 0.0728233, 0.0217709, -0.0383419, 0.1296900, 0.0720792, -0.0002758, 0.0869950, 0.1339810, 0.1771920, -0.0641624, -0.2432310, -0.5090030, -0.6462850, -0.3856790, -0.1861360, -0.0872939, -0.0215227, -0.0079253, -0.0071762, -0.0077304, -0.0022748, 0.0001757, 0.0004636, 0.0002562, 0.0012354, -0.0093115, -0.0188440, -0.0078165, -0.0382975, 0.0053321, -0.1098470, -0.1335190, -0.0967593, 0.0395086, 0.0659783, -0.0610230, -0.1293260, -0.1762520, -0.5777800, -0.5844370, -0.4288580, -0.3041000, -0.1356410, -0.1054620, -0.0277775, -0.0367365, 0.0036672, -0.0076362, -0.0062262, -0.0000176, -0.0004581, 0.0001400, 0.0039448, 0.0197126, 0.0661912, 0.2323610, 0.1613970, 0.1392790, 0.1627480, -0.0189697, 0.1808900, 0.0530323, 0.2090690, 0.0932897, 0.0769679, -0.0810485, -0.4028830, -0.4501940, -0.4208640, -0.2622330, -0.1665930, -0.1894550, -0.1192270, -0.0306179, -0.0062552, -0.0079740, -0.0013137, -0.0002676, -0.0004113, -0.0001796, 0.0001443, 0.0027101, 0.0380178, 0.0923027, 0.0851851, 0.1195410, 0.2461860, 0.2833790, 0.0766458, 0.0325695, 0.1307470, 0.2063850, 0.0850007, -0.0858265, -0.1137530, -0.2135270, -0.2019170, -0.1082110, -0.0698638, -0.0322386, 0.0012942, -0.0065671, -0.0023939, -0.0008322, -0.0011299, -0.0003631, -0.0003712, -0.0003341, -0.0002613, 0.0003114, -0.0002601, 0.0091853, 0.0441857, 0.0785105, 0.0890266, 0.1390410, 0.1214110, 0.1789940, 0.1593280, 0.2249160, 0.2119950, 0.1189720, 0.0375600, 0.0017869, 0.0275453, 0.0170713, 0.0022804, 0.0039419, 0.0061785, -0.0010427, 0.0000318, -0.0000101, -0.0001521, 0.0005248, -0.0009239, 0.0003836, -0.0002144, -0.0002982, 0.0002934, -0.0006532, 0.0039455, 0.0191656, 0.0168321, 0.0024106, 0.0080776, 0.0057343, 0.0053138, -0.0039337, 0.0333090, 0.0096618, 0.0065617, 0.0095448, 0.0284432, 0.0018409, 0.0003654, 0.0012231, 0.0039646, 0.0003290, -0.0003470, -0.0002399, -0.0002014, 0.0001640, -0.0007066, 0.0001878, 0.0001781, -0.0001053, -0.0003886, -0.0002616, -0.0005062, -0.0005816, 0.0000362, 0.0002207, 0.0003250, 0.0004926, -0.0003421, -0.0007278, 0.0001700, -0.0004090, 0.0005564, -0.0000475, -0.0000435, -0.0004103, -0.0005314, -0.0003147, -0.0008800, 0.0004864, 0.0000641, 0.0000023, 0.0002309, -0.0007615, 0.0002099, -0.0005068, -0.0001642, -0.0005044, -0.0003498, -0.0004657, -0.0006023, -0.0013852, -0.0043297, -0.0034118, -0.0107479, -0.0103300, -0.0164846, -0.0261771, -0.0148594, -0.0125921, -0.0191536, -0.0138407, -0.0101593, -0.0154565, -0.0249597, -0.0096902, -0.0026899, -0.0008217, 0.0002758, 0.0002166, -0.0001142, 0.0001204, 0.0002283, 0.0001243, 0.0000401, 0.0003388, -0.0019356, -0.0007567, -0.0032674, -0.0081871, -0.0132180, 0.0093207, -0.0021292, -0.0488547, -0.0408094, -0.0238968, -0.0890838, -0.0766542, -0.1173970, -0.1639330, -0.1483850, -0.1094830, -0.0787463, -0.0567282, -0.0205074, -0.0044174, 0.0073355, 0.0061776, 0.0000724, -0.0005498, 0.0002082, 0.0001161, 0.0050265, -0.0000887, -0.0022995, 0.0243547, 0.0097781, 0.0169161, 0.0208623, -0.0549161, -0.0575274, 0.0465681, 0.1438070, 0.1108860, -0.1486920, -0.1414960, -0.1714670, -0.3341680, -0.3640020, -0.2723300, -0.1882810, -0.1328850, -0.0534103, -0.0164193, 0.0001228, 0.0012326, -0.0045641, -0.0003942, 0.0002099, -0.0004327, 0.0142619, 0.0041851, 0.0057807, 0.1159730, 0.1696950, 0.1200670, 0.2177880, 0.0478740, 0.1268400, 0.0775592, 0.1267580, 0.0625014, -0.0453947, 0.0106894, -0.1445510, -0.3154090, -0.2842740, -0.3796680, -0.3429860, -0.2329670, -0.1260100, -0.0895413, -0.0596229, -0.0211336, -0.0026709, 0.0003162, 0.0004185, 0.0001815, 0.0026642, 0.0202133, 0.0938610, 0.2080350, 0.2278590, 0.1970210, 0.1471060, 0.0927077, -0.0836438, 0.0308996, 0.2900310, 0.1189230, 0.0487551, 0.1594970, 0.0325350, -0.0951297, -0.2171900, -0.5155130, -0.6563120, -0.4234280, -0.1991480, -0.1591460, -0.0619745, -0.0183972, -0.0049914, -0.0016176, 0.0000100, -0.0001699, 0.0021232, 0.0769029, 0.1797470, 0.1454550, 0.2269510, 0.1156070, -0.1038250, 0.0598274, 0.0202623, 0.0675251, -0.0188549, 0.1762570, 0.0764613, -0.0425260, 0.0978502, -0.0742053, -0.0171886, -0.3676770, -0.3737700, -0.3661760, -0.3023720, -0.1575550, -0.0686033, -0.0354096, -0.0147910, -0.0054960, -0.0003485, 0.0050998, 0.0005606, 0.1387010, 0.2618060, 0.0564988, 0.1077740, 0.0434373, -0.1040940, -0.0634260, 0.0151093, -0.0206121, -0.1561010, 0.1233920, 0.0490104, 0.1167740, 0.0263441, -0.1123130, -0.1265820, -0.2071110, -0.4399230, -0.5579820, -0.4242900, -0.2397920, -0.1552060, -0.0354514, -0.0091113, -0.0009117, -0.0003721, 0.0014476, 0.0039622, 0.0438888, 0.2508390, 0.0082545, -0.0828309, -0.1082400, -0.2777830, -0.1117400, 0.3038790, -0.2140120, 0.0681528, 0.2399080, 0.1324390, 0.1451940, 0.1813910, 0.1212890, -0.0250379, -0.1944800, -0.6497980, -0.6414770, -0.3904490, -0.2367780, -0.1703610, -0.0482952, -0.0020202, -0.0037291, 0.0000250, 0.0021696, 0.0052166, 0.0330731, 0.1593100, 0.1458190, -0.0031047, -0.1192940, -0.2772970, -0.1101070, -0.2028640, -0.1596710, 0.2854570, 0.2407510, 0.3696650, 0.5816680, 0.6006470, 0.1969810, -0.2672140, -0.4279400, -0.7105010, -0.5364120, -0.2862940, -0.1200300, -0.0537666, -0.0223378, -0.0050641, 0.0072600, 0.0000602, 0.0019560, 0.0063499, 0.0355754, 0.0537454, 0.1084130, 0.0137019, -0.1706000, -0.4330400, -0.3066030, -0.0481525, 0.0531931, -0.0062665, 0.2241220, 0.4519930, 0.5315640, 0.5945810, 0.1478620, -0.3050620, -0.4375080, -0.4895800, -0.3959160, -0.0941555, -0.0046896, -0.0828901, -0.0548064, -0.0028353, 0.0071373, 0.0002295, 0.0041363, 0.0128936, 0.0671394, 0.0655586, -0.0203770, -0.0499043, -0.1985530, -0.0454129, 0.0125162, -0.0180857, 0.3283770, 0.2865200, 0.3544880, 0.4444490, 0.3562590, 0.0408356, -0.4804030, -0.6821840, -0.5035640, -0.3109240, -0.2394140, 0.0479768, 0.1080470, -0.0302356, -0.0435688, -0.0071697, 0.0021626, -0.0002162, 0.0027640, 0.0075768, 0.0030059, -0.0229441, -0.0001393, -0.2001730, -0.2023790, -0.1424840, 0.0139318, 0.0813351, 0.0226751, 0.0438079, 0.0834424, 0.3932460, 0.2452920, -0.0197894, -0.3721670, -0.2797350, -0.2225900, -0.1343140, 0.0312103, 0.1825740, 0.1669360, 0.1345510, 0.1049960, -0.0060047, 0.0099861, 0.0008652, 0.0008288, 0.0024115, -0.0179065, -0.0688598, -0.1150300, -0.1341950, -0.1432630, -0.2070340, -0.1170400, -0.0615721, 0.1199440, 0.0141827, 0.1215990, 0.2562730, 0.1800720, 0.1156560, -0.1519250, 0.0450205, -0.0110277, 0.0734471, 0.0860318, 0.0970314, 0.0889713, 0.1528310, 0.1481980, 0.0573946, 0.0172386, -0.0008912, -0.0000021, 0.0003821, -0.0118698, -0.0623290, -0.0685107, -0.1038750, -0.2041460, -0.1071280, -0.1346340, -0.0675979, -0.0665138, -0.1162950, 0.0142157, 0.1022410, 0.1298410, -0.1323390, -0.2727790, -0.1551050, 0.1266250, 0.0929832, 0.2292540, 0.0688824, 0.0454903, -0.0117393, 0.1228660, 0.0546403, 0.0010215, -0.0003924, -0.0004034, 0.0003221, 0.0338098, -0.0874360, -0.0757154, 0.0270597, 0.0858976, 0.2303320, -0.0181092, -0.0632188, -0.0277747, -0.1428640, 0.1797530, 0.1672290, 0.2272780, -0.0407641, -0.0071199, -0.1403850, 0.0657331, 0.2053140, 0.1258630, 0.2758300, 0.1012100, 0.0833045, 0.0576493, 0.0897147, 0.0115630, 0.0003604, 0.0004986, -0.0004543, 0.0260027, -0.0617183, -0.1136530, 0.0541767, 0.3259960, 0.1953430, 0.2918990, -0.0155198, -0.1435190, -0.1061180, -0.0170525, 0.2526370, -0.0268704, -0.2008290, -0.2117790, 0.0714046, -0.0187616, -0.0013667, 0.0253697, 0.1350000, 0.1422060, 0.1768780, 0.0402485, 0.1244040, 0.0242898, -0.0000558, -0.0000472, 0.0006448, -0.0154115, -0.0711613, -0.1725450, 0.0195381, 0.1106220, -0.0873376, -0.0227855, -0.1684040, -0.2160890, -0.1557340, -0.0283050, 0.1239570, -0.1590810, -0.1127290, -0.0163808, -0.0139170, 0.0508679, -0.0101584, 0.1488100, 0.1564930, 0.1128630, 0.1665500, 0.0857429, 0.0462664, 0.0061601, 0.0016705, 0.0003365, -0.0002011, -0.0179314, -0.0220794, -0.0941638, -0.0655182, -0.1993970, -0.1027800, -0.0312848, 0.0977680, 0.0117110, -0.1496190, -0.0669796, -0.2234640, -0.1545460, -0.0623073, 0.0589438, 0.0285173, 0.1561030, 0.1319780, 0.1229940, 0.2698920, 0.1940330, 0.1534000, 0.0794330, 0.0105782, 0.0058137, 0.0000995, -0.0022271, -0.0581662, -0.0703254, -0.0069122, -0.0515867, -0.3143860, -0.1659190, -0.1319790, -0.0510441, 0.0029781, -0.1886610, -0.1806860, -0.0301084, 0.0460746, -0.1134940, 0.0554554, 0.0540202, 0.0821923, 0.1341280, 0.1999690, 0.0162622, 0.1443060, 0.0940426, 0.0250580, 0.0473722, 0.0281785, 0.0016112, 0.0002284, -0.0053676, -0.0496818, -0.0628296, -0.0861603, -0.1258000, -0.0736600, 0.0766817, 0.0616148, 0.1343790, -0.0500499, -0.1097640, -0.1247700, -0.0643484, 0.0007026, -0.2889970, -0.0716935, -0.1275010, 0.0125131, -0.0673526, 0.0588380, -0.0345651, -0.0527153, 0.0281442, -0.0569541, -0.0630114, 0.0079139, -0.0003358, 0.0000671, 0.0003586, 0.0052504, 0.0029209, -0.0910388, -0.1887040, -0.1519330, -0.1502980, -0.1044120, -0.0676384, -0.0908218, -0.0547860, -0.1012660, -0.2866530, -0.0755560, -0.0474645, 0.0304731, -0.1347440, -0.0761485, -0.0288124, -0.1766800, -0.1723190, -0.0607643, -0.0557320, -0.1358480, -0.0718046, -0.0002833, -0.0000091, -0.0003117, -0.0003556, 0.0034803, 0.0172027, 0.0155366, -0.1048760, 0.0035633, -0.1029860, -0.1571740, -0.1552900, -0.0153199, -0.1870220, -0.1527220, -0.0541923, -0.1970850, -0.1225000, -0.2421660, -0.1914780, 0.0674154, 0.0339835, 0.0663204, 0.0421276, 0.0018587, -0.1486480, -0.1382050, -0.0699673, -0.0086210, 0.0002301, 0.0001539, 0.0002668, 0.0031386, 0.0157671, 0.0271898, -0.0338912, -0.0853320, -0.0171999, -0.0667554, 0.0357815, -0.0013014, 0.0732599, -0.1249300, 0.0901337, -0.2486330, -0.0562081, -0.2112980, 0.0233428, -0.0440982, -0.1513900, 0.0655051, -0.0000644, -0.0635499, -0.1544310, -0.1218790, -0.0460691, -0.0045075, -0.0003013, 0.0000678, 0.0002163, 0.0014475, 0.0073728, 0.0532493, 0.0549506, 0.0726748, 0.0601501, 0.0569359, 0.0051788, -0.1076660, -0.0204428, -0.2680650, -0.0139870, 0.1203740, -0.1801760, -0.1451660, -0.0614430, -0.1899900, -0.1293680, -0.1366270, -0.0093541, -0.0509404, -0.1350600, -0.0592204, 0.0083264, 0.0012764, -0.0005647, -0.0000061, 0.0002617, -0.0003814, -0.0009081, 0.0507800, 0.1091200, 0.1363290, 0.1611610, 0.1386020, 0.0884276, 0.1068240, -0.0143849, -0.0006756, 0.1589810, 0.1170970, -0.0740734, -0.0683241, -0.0057572, -0.0231747, -0.1248440, -0.0724567, -0.0616222, -0.0426889, -0.0885698, -0.0460985, 0.0008707, 0.0012552, 0.0001483, -0.0007646, 0.0005628, 0.0000153, 0.0002049, -0.0004326, -0.0017847, 0.0012498, 0.0031898, -0.0090481, -0.0103659, -0.0194215, -0.0398625, -0.0986267, -0.0273553, -0.0145461, -0.0394664, -0.0571435, -0.0084161, 0.0142273, -0.0281878, -0.0338712, -0.0086519, 0.0028343, -0.0010377, -0.0001125, 0.0004485, -0.0002100, -0.0000868, -0.0001643, 0.0001040, 0.0004305, -0.0000480, 0.0000347, 0.0002917, -0.0014350, -0.0069379, -0.0062428, 0.0005399, 0.0022842, 0.0095359, 0.0089734, 0.0215562, 0.0110654, 0.0009271, -0.0038093, 0.0035131, -0.0059083, -0.0021360, 0.0002932, 0.0211138, 0.0115684, 0.0005104, -0.0000301, -0.0002339, 0.0000056, 0.0000281, 0.0000295, 0.0002183, -0.0000558, 0.0004106, 0.0002828, 0.0004565, 0.0005312, -0.0007773, 0.0002524, -0.0000439, 0.0003163, 0.0003222, 0.0000624, -0.0001572, 0.0003484, -0.0000793, -0.0000579, -0.0003269, 0.0001572, -0.0003921, 0.0000623, -0.0003408, -0.0004286, -0.0006317, 0.0002031, 0.0000778, 0.0000157, -0.0005066, -0.0005434, 0.0005513, -0.0001165, 0.0000911, -0.0006849, -0.0001370, 0.0007609, 0.0020404, 0.0079116, 0.0023406, 0.0034690, 0.0096038, 0.0059545, 0.0037658, -0.0071101, -0.0074269, 0.0264595, 0.0119700, -0.0010317, -0.0006454, -0.0019989, -0.0012257, 0.0001659, -0.0002405, -0.0000841, 0.0005202, -0.0001839, 0.0003484, 0.0001432, 0.0001538, 0.0004567, 0.0009075, 0.0002574, 0.0008248, 0.0008550, 0.0036607, 0.0088053, 0.0129552, 0.0320688, 0.0335594, 0.0417600, 0.0200626, -0.0093168, -0.0879581, -0.1041070, -0.0919848, -0.0658896, -0.0845701, -0.0353545, -0.0152558, -0.0077455, 0.0004555, 0.0003541, 0.0000668, -0.0003590, 0.0004574, -0.0001660, 0.0003305, -0.0015141, 0.0027863, 0.0030113, -0.0123608, -0.0128392, -0.0637970, -0.0559547, 0.0601845, -0.0010865, 0.0098700, 0.0163136, 0.0009310, -0.0946305, -0.2576070, -0.1961970, -0.1441410, -0.2020680, -0.1713680, -0.1817240, -0.0628933, -0.0183009, -0.0064457, -0.0012606, -0.0001295, -0.0002644, -0.0001085, 0.0000146, -0.0005231, -0.0061676, -0.0035635, -0.0027339, -0.0463181, -0.0356403, -0.0398224, -0.0877511, 0.0357038, -0.0737299, 0.0247754, 0.1338820, -0.0263211, 0.0027766, -0.1147440, -0.0789612, 0.1150840, -0.1261200, -0.2012950, -0.0636739, -0.1145070, -0.0470784, 0.0216345, -0.0013528, -0.0037582, 0.0013086, 0.0007230, -0.0003197, 0.0001836, -0.0017397, -0.0108787, -0.0331719, -0.1033160, -0.0257253, -0.1042720, 0.0010404, -0.0565232, 0.1291920, 0.2984990, -0.0390513, -0.1569860, -0.2742410, -0.1912930, -0.1203440, -0.0148796, 0.0737500, -0.0026340, 0.1007890, 0.1003030, -0.0198224, -0.1004220, -0.0097532, 0.0153389, 0.0086618, -0.0001673, 0.0004347, -0.0003852, -0.0102386, -0.0450347, -0.1040700, -0.2003480, -0.2196080, -0.0889848, 0.1398290, 0.1119560, 0.0564116, 0.2266090, -0.0417047, -0.1237130, 0.0159865, 0.0146978, 0.1052320, 0.1940820, 0.1232660, 0.0050087, 0.0411575, 0.0928276, 0.0377355, -0.0535539, -0.0929458, -0.0010918, -0.0006128, -0.0009180, 0.0000864, -0.0118333, -0.0002285, -0.0781401, -0.1167500, -0.0946534, -0.1069220, -0.1169820, 0.1744830, 0.2788830, 0.3583500, 0.0484169, -0.1626050, -0.1305810, -0.0664700, 0.0729263, 0.1205790, 0.1504130, 0.1153920, -0.1276520, 0.0007176, 0.0900260, 0.0847215, -0.1031600, -0.0461237, 0.0240484, -0.0013357, -0.0001288, 0.0049834, -0.0078103, -0.0052089, -0.0513886, -0.1119870, -0.1130460, 0.0186977, -0.0864195, 0.2555340, 0.2449560, 0.2172080, 0.0221959, -0.3546430, -0.2890300, -0.0331841, 0.0546609, 0.3003640, 0.1521140, 0.0133040, -0.1592830, -0.1693280, -0.0307541, -0.1571880, -0.0173387, 0.0206741, 0.0028404, 0.0017213, -0.0001018, -0.0003399, -0.0094122, -0.0164129, -0.0273560, -0.0785674, -0.0289385, -0.0512530, -0.1154490, 0.0094638, 0.0987883, 0.4158780, 0.0400306, -0.1684230, -0.3886300, -0.3088270, 0.1553880, 0.0819179, -0.0448294, -0.0187283, -0.0845771, -0.1109580, -0.1121550, -0.2207290, -0.0470901, 0.0598748, -0.0158578, 0.0035826, -0.0020666, -0.0003899, -0.0073253, -0.0141058, -0.0310005, 0.0463911, 0.0048069, 0.0624792, -0.0140530, 0.1944480, 0.2229570, 0.2395870, 0.2493090, -0.1007320, -0.4282590, 0.1112600, 0.1727860, 0.1020450, -0.0990000, -0.0319403, -0.1579420, -0.1449980, 0.0018431, -0.0983559, 0.0999668, 0.1344090, -0.0045574, 0.0030061, -0.0013793, 0.0001980, -0.0058971, -0.0395523, -0.0579685, -0.0397618, -0.1037470, -0.0133587, 0.1552480, 0.2226410, 0.2092560, 0.2925720, 0.3274330, 0.0096979, -0.1689840, 0.0849865, 0.0205451, 0.1944840, 0.0834363, -0.1572610, -0.0467848, 0.1084860, 0.3016870, 0.1354730, 0.1698720, 0.2036270, 0.0341623, 0.0022124, -0.0003014, 0.0008087, -0.0040835, -0.0344034, 0.0322447, 0.1061100, -0.0140870, 0.0405475, 0.0274406, 0.1162760, 0.1337380, 0.1823610, 0.1891600, -0.1688440, -0.1639760, -0.2581270, -0.3001670, -0.0781090, 0.0108940, -0.3547570, 0.0540011, 0.0426588, 0.2289590, 0.1305280, 0.2699830, 0.2015140, 0.0352032, 0.0037124, -0.0009930, 0.0000809, -0.0017513, -0.0285764, 0.0136483, 0.1221100, 0.1051840, 0.0031863, 0.3064850, 0.1485150, 0.1150110, 0.2553720, 0.1022980, 0.1187980, -0.0969626, -0.0224238, -0.0233579, -0.0198118, -0.0749393, -0.3826790, 0.0383166, 0.0781083, 0.2143840, 0.3870280, 0.3035150, 0.1241720, 0.0519732, 0.0120805, 0.0008711, 0.0002619, -0.0028045, -0.0177328, -0.0128121, 0.0494628, 0.0477726, 0.1732720, 0.3547990, 0.0574153, 0.0812478, 0.3482720, 0.4087990, 0.1568810, 0.1710750, -0.0990173, -0.1992260, 0.0706070, -0.0427238, 0.0203041, -0.0771414, 0.0961845, 0.0877210, 0.2346010, 0.0298703, 0.0000207, 0.0729084, 0.0255485, 0.0001343, 0.0000963, -0.0031458, -0.0015209, -0.0120515, 0.0653807, -0.0285733, -0.0187823, 0.1133910, -0.0058369, 0.2283310, 0.3665830, 0.4092470, 0.2738000, 0.0665765, -0.0853479, -0.3276880, -0.1024200, -0.0991701, -0.1253470, -0.3766660, -0.3316690, -0.3308740, -0.0951478, -0.0524637, -0.0253852, 0.0914106, 0.0145696, 0.0019945, 0.0007319, -0.0010271, 0.0013600, -0.0578402, 0.0632469, 0.0030939, 0.0662616, -0.0583708, 0.0614370, 0.1691520, 0.2770470, 0.2899250, 0.2651690, -0.0459692, -0.0365816, -0.2201440, 0.0296890, -0.1166890, -0.1872980, -0.5289610, -0.3124390, -0.3962160, -0.1163030, -0.0944552, -0.0782447, 0.1279290, 0.0374148, 0.0085507, -0.0005438, -0.0005732, -0.0143951, -0.0104017, 0.0029266, -0.0625344, 0.0402394, -0.0717680, 0.1289750, 0.3543940, 0.3529780, 0.1444690, 0.2018820, -0.0938426, -0.1549140, -0.1217950, -0.1309730, -0.1685370, -0.1685320, -0.4199290, -0.0928374, -0.3840090, -0.1658800, -0.1907300, 0.0293117, 0.1744970, 0.0398375, 0.0281946, 0.0001907, -0.0006072, -0.0245564, -0.0874283, -0.0274773, -0.0668447, -0.0066311, -0.0489734, 0.0245550, 0.1847890, 0.3634870, 0.1712900, 0.1220280, -0.1599720, -0.1750590, -0.3329650, -0.2796440, -0.2512240, -0.2046730, -0.1813160, -0.1400900, -0.2553530, -0.1304810, -0.1716930, 0.0779747, 0.0787566, 0.0041880, 0.0012629, 0.0000700, -0.0013308, -0.0229680, -0.1624950, -0.0281636, -0.0295145, -0.0173867, 0.1343510, 0.0811121, 0.1056260, 0.2316970, 0.1304990, 0.2399420, -0.0239421, -0.2750690, -0.0978829, -0.2205320, -0.3258760, -0.1255320, -0.0761698, -0.1765630, -0.1423460, 0.0064975, 0.0704877, 0.0647823, 0.0195891, 0.0074745, -0.0002377, -0.0008508, 0.0001267, -0.0050446, -0.0962265, -0.0319806, 0.0783127, -0.0170637, 0.0299457, 0.0083824, -0.0349684, 0.1811860, 0.1785260, 0.2161070, -0.0794235, -0.2551300, -0.0850724, -0.1810570, -0.1609730, -0.2411210, -0.0648444, -0.2371070, -0.1332220, 0.0660449, 0.1258060, 0.1195590, 0.0442293, 0.0017224, 0.0004019, -0.0004732, -0.0004541, 0.0148303, -0.0074055, -0.0402029, 0.0499997, -0.0348202, -0.0187718, -0.0071483, 0.2018630, 0.0535898, -0.0205136, -0.0730105, 0.0764103, -0.1041210, -0.0247748, -0.0658513, 0.0397326, -0.2119040, -0.1304170, -0.0542134, 0.2220270, 0.2500110, 0.2341590, 0.1029810, 0.0196146, 0.0048304, -0.0000085, 0.0011103, -0.0003370, -0.0025846, 0.0344332, -0.0680921, -0.1615430, -0.0330722, 0.0521257, 0.1383710, 0.1587520, 0.0521066, 0.0216594, 0.0025500, 0.1483870, 0.0619691, -0.2336740, -0.0372527, -0.0932098, -0.0921590, -0.2741280, 0.0953425, 0.1723650, 0.1536800, 0.1881080, 0.0656563, 0.0168642, -0.0015684, 0.0003779, -0.0001555, -0.0001108, -0.0115213, -0.0338696, -0.1623250, -0.1490490, -0.1242540, -0.2130310, 0.1212600, -0.0562345, -0.1019800, -0.1006660, 0.0618265, 0.1311580, -0.0062381, -0.1701140, 0.1471560, 0.1699170, 0.0050884, -0.0716602, 0.1034060, 0.1901140, 0.2203800, 0.1686470, 0.0434051, 0.0057365, -0.0022663, 0.0004397, 0.0000092, -0.0003192, -0.0044332, -0.0568887, -0.1287550, -0.1782850, -0.2693350, -0.3148260, -0.2507870, -0.1620750, -0.1922610, -0.2037510, 0.0895781, -0.1212280, -0.3719100, -0.0686268, 0.0866433, 0.0419651, 0.0615240, 0.0888305, 0.1615460, 0.0982391, 0.1204820, 0.0915323, 0.0412418, 0.0053963, 0.0004682, -0.0001905, -0.0004664, 0.0006800, -0.0000517, -0.0027667, -0.0300787, -0.0791827, -0.1430470, -0.2007430, -0.3089770, -0.2396280, -0.2206720, -0.1780270, -0.3837670, -0.0845504, 0.0232637, 0.0653252, 0.0619929, -0.0444092, -0.0690681, 0.0138388, 0.1047620, 0.0831985, 0.0368474, 0.0158498, 0.0034490, -0.0003308, -0.0000920, -0.0002522, 0.0002173, -0.0005196, -0.0006158, 0.0001833, 0.0047201, 0.0146943, 0.0032298, -0.0094971, -0.0387807, -0.0943111, -0.1574580, -0.1246740, -0.0208098, -0.0561644, 0.0201696, -0.0550226, -0.0398824, -0.0185892, 0.0217627, 0.0058527, 0.0569228, 0.0702278, 0.0257450, 0.0037439, -0.0002534, -0.0001490, -0.0000731, 0.0005155, 0.0001138, -0.0001907, -0.0003781, -0.0004038, -0.0005246, -0.0023181, -0.0014885, 0.0072994, 0.0047515, -0.0050924, -0.0075615, -0.0008953, -0.0061507, -0.0305698, -0.0104453, 0.0059671, -0.0089714, -0.0167499, 0.0102800, 0.0226519, 0.0117369, 0.0075996, 0.0128401, -0.0010943, -0.0006304, 0.0001409, 0.0005462, -0.0003452, -0.0002502, 0.0000362, 0.0000295, 0.0002819, 0.0000876, -0.0000799, 0.0000073, 0.0007902, 0.0004071, 0.0004051, 0.0002302, -0.0000207, -0.0017000, -0.0026239, -0.0000710, -0.0000815, -0.0001808, 0.0001667, 0.0000087, 0.0002043, -0.0002497, -0.0004065, 0.0003413, 0.0002366, 0.0001323, -0.0000760, 0.0000420, -0.0001107, 0.0002143, 0.0005245, -0.0002535, 0.0001718, -0.0005747, -0.0002220, -0.0137931, -0.0230482, -0.0395069, -0.0133871, -0.0246557, -0.0269497, -0.0426819, -0.0455568, -0.0058629, -0.0086601, -0.0177005, -0.0221096, -0.0232584, -0.0255156, -0.0232240, -0.0089347, -0.0052979, -0.0036917, 0.0008983, -0.0004325, 0.0001107, 0.0003928, 0.0004302, 0.0001331, -0.0001006, -0.0017864, -0.0020007, -0.0004617, -0.0136754, -0.0499909, -0.0689179, -0.0568514, -0.0744141, -0.1141110, -0.1663320, -0.1377200, -0.1233130, -0.1016740, -0.0833990, -0.0539130, -0.0478736, -0.0690102, -0.0702381, -0.0635057, -0.0286966, -0.0290688, -0.0188371, -0.0045347, 0.0003803, -0.0002497, -0.0001229, -0.0001695, 0.0000321, -0.0039863, -0.0070009, -0.0162604, -0.0835262, -0.1286840, -0.1803820, -0.2310710, -0.1995600, -0.2441830, -0.2684890, -0.2912020, -0.1893860, -0.1354280, -0.1236280, -0.0687654, -0.0128935, -0.0622408, -0.1476440, -0.0780961, -0.0083899, -0.0861224, -0.0748490, -0.0018250, -0.0090238, 0.0001006, 0.0000007, 0.0002811, 0.0015358, 0.0009048, -0.0176935, -0.0523060, -0.1092250, -0.1565410, -0.3426220, -0.4830070, -0.4255350, -0.2562640, -0.2969180, -0.4678820, -0.4717540, -0.3750350, -0.3500110, -0.1407680, -0.1471870, -0.2057560, -0.1580010, 0.0681431, 0.0480061, 0.0110870, 0.0466276, 0.0268669, 0.0165335, -0.0022379, 0.0000889, 0.0002453, -0.0019257, -0.0026059, -0.0703177, 0.0168345, -0.0848984, -0.1224890, -0.0970378, -0.3129180, -0.4865020, -0.2032230, 0.1018630, -0.2596230, -0.2692480, -0.4252300, -0.2917970, -0.3042270, -0.4021080, -0.4091890, -0.1707020, -0.0917971, 0.0126353, -0.0117673, 0.0473948, 0.0703800, 0.0037137, 0.0006856, 0.0000901, -0.0000441, 0.0094084, 0.0342886, -0.0082329, 0.1325330, -0.0328127, -0.0720505, -0.0507725, 0.1189190, 0.1153840, -0.1051710, 0.1714070, 0.0765178, 0.0932844, 0.0846039, 0.0441393, 0.1369360, 0.0253561, 0.1046180, 0.0442129, 0.0677383, -0.0761519, -0.0257728, 0.0607607, 0.0950142, 0.0623405, -0.0010878, 0.0001019, 0.0030618, 0.0304799, 0.0860009, -0.0419873, -0.0521844, 0.0835789, 0.0523714, 0.1890050, 0.1887380, 0.0236923, -0.0196388, 0.1016320, 0.1685760, 0.0597066, 0.1283710, 0.4340450, 0.1868930, -0.0364375, 0.1601090, 0.1452870, 0.0537966, -0.0147880, 0.0123823, 0.0945468, 0.1003720, 0.0551693, -0.0034192, -0.0061744, 0.0047282, 0.0189724, 0.0622086, -0.0337063, -0.0110919, 0.0877731, 0.0431403, 0.2569930, 0.1679450, 0.1286500, 0.2149230, 0.0183661, -0.1947960, 0.0336064, 0.1954450, 0.1896220, -0.0130768, 0.1415690, 0.0204401, 0.0201782, 0.1644050, 0.1499710, 0.2150620, 0.2748450, 0.1923710, 0.0290243, 0.0045200, 0.0003936, 0.0058647, 0.0027616, 0.0575943, 0.0158164, -0.0699857, 0.0607892, 0.0228079, 0.2214270, 0.1352270, 0.0707580, 0.2242600, 0.1344000, -0.0297253, -0.0718346, 0.0396558, 0.0926580, 0.2023960, 0.0264977, -0.0411041, -0.0355175, 0.2265840, 0.2526320, 0.2233830, 0.1091800, 0.1925390, 0.0861878, 0.0701819, 0.0005058, 0.0017620, -0.0108119, 0.0241469, 0.0750974, 0.0316776, 0.1057570, 0.1495670, 0.2040790, 0.1475850, 0.0934920, -0.0689586, -0.0855132, -0.0754873, -0.2306790, 0.0589702, -0.0268368, -0.1023190, 0.1228140, 0.1677260, 0.0836287, 0.1207210, 0.1324330, 0.0123082, 0.0780717, 0.1717730, 0.0676904, 0.0235807, 0.0004505, 0.0026330, 0.0158686, 0.0193548, 0.1124260, 0.1276190, 0.1790670, 0.1568930, 0.3389780, 0.3812660, 0.2472370, 0.1395960, 0.1280930, 0.0888431, -0.0672034, -0.0552276, -0.1227260, -0.0371088, -0.1610900, -0.1306320, -0.1364800, -0.0548103, 0.0586123, -0.0996825, -0.0624050, 0.0461957, 0.0398012, 0.0070181, 0.0002808, 0.0041657, 0.0341889, 0.0493705, 0.1505570, 0.2275190, 0.2497710, 0.1023410, 0.2767220, 0.2884000, 0.2770410, 0.2010990, 0.1327360, 0.0732045, -0.3327220, 0.0470542, -0.0104065, 0.0436066, 0.1049010, 0.0357382, -0.1032220, -0.0478630, -0.0999666, -0.2369020, -0.2279990, 0.0902398, 0.0899203, 0.0192232, -0.0001312, 0.0012980, 0.0206843, 0.0011072, 0.1570430, 0.2543740, 0.2726730, 0.2676800, 0.1440430, 0.3101280, 0.4164390, 0.4723910, 0.1014840, -0.0112794, -0.2471230, 0.1996920, 0.0886837, 0.1593990, -0.0306247, -0.0508491, -0.0293457, -0.0160305, -0.0555561, -0.2308010, -0.1551260, 0.0573367, 0.0328077, -0.0032107, -0.0001349, 0.0007290, 0.0048594, -0.0275669, 0.1175360, 0.1023910, 0.0913094, 0.1615660, 0.2273840, 0.1715350, 0.1738050, 0.1863930, 0.3339100, -0.0180003, -0.0303182, 0.2136390, 0.2966330, 0.2440600, -0.0740015, 0.1405900, -0.0779730, -0.1023230, -0.1557060, -0.0982640, -0.1149310, -0.0308027, 0.0074037, -0.0003759, -0.0001023, -0.0002336, -0.0049854, 0.0061180, 0.0357135, -0.0782326, 0.1502150, -0.0334536, 0.1004180, -0.0283805, 0.1261230, 0.2496820, 0.1809050, -0.0598907, 0.0351912, 0.3020050, 0.1918220, 0.3557550, -0.0308803, -0.1106070, -0.0923401, 0.0890671, 0.0083099, -0.1453340, -0.2155450, -0.0558153, 0.0381532, 0.0016285, -0.0000111, -0.0002387, -0.0083993, 0.0147330, 0.0172359, -0.2020190, -0.0138001, 0.0069473, 0.0281861, 0.0496227, -0.0782163, -0.0282977, 0.1691810, 0.3817520, -0.0184114, 0.2049450, 0.2507550, 0.3298620, -0.0923637, -0.1986110, -0.0737086, 0.0843360, -0.0010876, -0.1406800, -0.2249350, -0.0449951, 0.0382457, 0.0073525, 0.0003622, 0.0003109, -0.0057067, -0.0307372, -0.0390344, -0.1291900, 0.0267986, 0.0486181, -0.0701311, 0.0241412, -0.2376750, -0.0419931, -0.0726837, 0.2930870, 0.1647850, 0.2274150, 0.1718110, 0.1960910, 0.2068820, -0.2118660, -0.2188440, -0.0481661, 0.0809509, -0.0983523, -0.0631993, -0.0669966, 0.0327398, -0.0190358, 0.0010673, 0.0002616, 0.0009723, -0.0946144, -0.1271880, -0.0007755, -0.0669581, 0.0569433, 0.0119458, -0.1438630, -0.0046970, 0.2269710, 0.0920179, 0.0205885, -0.0428112, -0.1966560, -0.1542640, 0.0300296, -0.0424651, -0.0267185, -0.0572565, -0.0745505, -0.0352740, -0.1806910, -0.1541450, -0.0492923, 0.0279936, -0.0029472, 0.0000899, 0.0046667, 0.0003608, -0.1256120, -0.2378710, -0.1744590, -0.2350190, -0.1530740, -0.0015704, -0.1027380, -0.1920770, -0.1960100, -0.2376460, -0.3446390, -0.4560620, -0.3005760, -0.0867196, -0.0428381, -0.1514440, 0.0574496, -0.0514687, -0.1774810, -0.3048150, -0.2135940, -0.0982747, -0.0207255, 0.0028213, -0.0013981, -0.0001297, -0.0024570, -0.0042903, -0.1435650, -0.3128800, -0.4003990, -0.4064360, -0.4182030, -0.3337530, -0.2821950, -0.2373260, -0.3273530, -0.3289720, -0.1100830, -0.2487770, -0.2247450, -0.1382010, -0.0667853, -0.3530380, 0.0287994, -0.0561031, -0.1188180, -0.1537990, -0.0877098, -0.0696500, -0.0209458, -0.0015222, 0.0005153, -0.0000494, -0.0000872, -0.0057328, -0.1636290, -0.1791640, -0.3229570, -0.4544240, -0.4497370, -0.3446870, -0.3416720, -0.3454260, -0.2737000, -0.0829352, -0.1943540, -0.2663780, -0.2395620, -0.2497190, -0.2552010, -0.2654210, 0.1044620, 0.1023040, 0.1359830, -0.1173200, -0.0606071, 0.0072847, -0.0107467, -0.0101387, -0.0003490, -0.0001332, -0.0003706, -0.0086164, -0.0856391, -0.1241710, -0.1934780, -0.2856550, -0.1199690, -0.2433940, -0.3028370, -0.1751360, -0.1173170, -0.0092995, -0.2610550, -0.1104650, -0.2482400, -0.1746900, -0.1874070, -0.2508720, 0.0383892, 0.0201130, 0.0018047, -0.0973292, -0.0099568, 0.0226763, -0.0015072, 0.0057002, 0.0001726, 0.0001742, -0.0002911, -0.0223926, -0.0428286, 0.0271626, -0.0012892, -0.0082612, 0.0811104, -0.1066690, -0.2983530, -0.1579390, -0.1642570, -0.2946990, -0.2250000, -0.0362273, -0.0252441, -0.0003170, -0.1966430, -0.1863110, -0.1105150, 0.0321144, 0.0352324, -0.0252548, -0.0122785, 0.0046517, 0.0083045, 0.0014199, -0.0003235, -0.0002222, -0.0004301, -0.0165599, -0.0124277, 0.0938631, 0.2090730, 0.1976900, 0.1535090, 0.0257744, -0.1157600, 0.1057500, 0.1857060, 0.0119044, -0.0546699, -0.0340467, -0.0155050, 0.0743478, 0.1129920, 0.0556265, 0.1405740, 0.1643180, 0.1411740, 0.0290626, -0.0063936, -0.0242097, -0.0116053, -0.0000244, -0.0003006, -0.0002937, -0.0003478, -0.0025773, 0.0123618, 0.0915796, 0.1054600, 0.1005030, 0.1678210, 0.1515950, 0.2299890, 0.2709810, 0.2448450, 0.2315380, 0.1572200, 0.2709910, 0.4021420, 0.3288980, 0.2619880, 0.1421230, 0.0825886, 0.1154740, 0.1226900, 0.0299560, 0.0086268, 0.0018982, -0.0002021, -0.0004450, -0.0000192, 0.0004893, -0.0002853, 0.0002532, -0.0006186, -0.0023488, -0.0241889, -0.0039923, 0.0474663, 0.0735478, 0.1247820, 0.0218181, -0.0139362, 0.1265220, 0.1405290, 0.1372890, 0.1232660, 0.0658677, 0.0831588, 0.0528409, 0.0267559, 0.0546051, 0.0512548, 0.0213156, 0.0009021, 0.0004290, -0.0003787, -0.0001958, 0.0004776, -0.0003825, 0.0002804, -0.0002858, -0.0004696, -0.0000881, 0.0005430, 0.0017944, 0.0016669, 0.0018064, 0.0082410, 0.0275984, 0.0112246, 0.0068803, 0.0075305, 0.0057478, 0.0107440, 0.0054974, 0.0058037, 0.0052493, 0.0086645, 0.0158176, 0.0125817, 0.0216688, 0.0050437, 0.0003639, 0.0002201, -0.0000933, -0.0002314, 0.0000976, -0.0001885, -0.0003011, -0.0003722, -0.0000573, 0.0004728, 0.0002422, -0.0002277, -0.0003020, 0.0003227, -0.0002514, -0.0004802, -0.0000188, -0.0000538, -0.0000304, 0.0001489, -0.0002186, 0.0002069, -0.0005853, 0.0001562, -0.0004783, 0.0000031, -0.0001169, -0.0002959, 0.0001845, -0.0005218, -0.0006790, -0.0004447, 0.0000444, -0.0000998, -0.0000054, -0.0001372, 0.0006902, 0.0007000, 0.0004619, 0.0023825, 0.0052010, 0.0037952, 0.0043856, 0.0030112, 0.0062304, 0.0100157, 0.0081807, 0.0075646, 0.0118290, 0.0084160, 0.0057329, 0.0052808, 0.0054389, 0.0033841, 0.0024706, 0.0024370, -0.0000143, 0.0004684, 0.0004156, 0.0002440, -0.0003581, 0.0000517, 0.0003866, 0.0000520, 0.0002292, -0.0005974, 0.0008114, 0.0029688, 0.0043389, 0.0069503, 0.0120080, 0.0282793, 0.0552654, 0.0882852, 0.0814983, 0.0527220, 0.0314680, 0.0188332, 0.0329948, 0.0661945, 0.0336009, 0.0171960, 0.0098381, 0.0035778, 0.0019381, 0.0008340, 0.0005024, -0.0005333, -0.0004456, -0.0001290, 0.0006486, -0.0002775, -0.0027476, 0.0224045, 0.0282552, 0.0442605, 0.0348613, -0.0192651, 0.0053959, 0.0798569, 0.0990396, 0.1765370, 0.1439590, 0.0173476, 0.0357597, 0.0206587, 0.0106911, -0.0254209, -0.0646583, -0.0815985, -0.0026993, 0.0146960, 0.0054487, 0.0012088, 0.0006230, 0.0001210, -0.0002576, -0.0001190, 0.0008808, 0.0014701, 0.0100933, 0.0580711, 0.0711618, 0.0221253, 0.1226850, 0.0763694, 0.2091470, 0.2448440, 0.1750150, 0.1010400, 0.0852238, 0.0745841, -0.0225100, -0.1535670, -0.1499560, -0.0080894, -0.0703908, -0.1165460, -0.0881302, -0.0656728, -0.0289094, 0.0049101, 0.0095529, 0.0013667, 0.0003141, -0.0003427, 0.0012880, 0.0137138, 0.0937785, 0.1590540, 0.1962010, 0.2230340, 0.2345030, 0.0794115, -0.0469380, -0.0244871, 0.1301820, 0.1833550, -0.0263169, 0.2205540, -0.1043350, -0.2461870, -0.2484440, -0.0319169, -0.0563723, -0.1244690, -0.2150310, -0.1760720, -0.0336256, 0.0177513, 0.0077884, -0.0004086, 0.0005398, 0.0003676, -0.0114427, 0.0499944, 0.1257000, 0.0302022, 0.1124890, 0.2469300, 0.2159160, 0.1319120, 0.0091022, -0.2017830, -0.0929717, -0.0515742, -0.1274690, 0.1777110, 0.4350630, 0.2399750, 0.0106940, -0.4079640, -0.1983950, -0.0478019, -0.3288840, -0.3349450, -0.1213020, 0.0113614, 0.0018096, 0.0014947, 0.0000699, 0.0020408, -0.0125670, 0.0806722, 0.1002060, -0.1234350, -0.0542490, 0.1089580, 0.0794114, -0.0629272, -0.1213490, -0.3286120, -0.1401370, -0.2677410, -0.1076900, 0.3840240, 0.1626630, 0.1269150, 0.0033532, -0.0491679, -0.0618313, -0.0991165, -0.3195300, -0.4046600, -0.2925820, -0.0704778, 0.0033343, 0.0006387, -0.0020104, 0.0009435, 0.0040170, 0.0629343, 0.0540399, -0.0313263, -0.0774119, -0.0029084, 0.0906627, 0.0728246, 0.1001860, -0.2961250, -0.3176760, -0.1605650, 0.0995559, 0.2491170, 0.3339820, -0.0118565, 0.1935990, 0.1491380, 0.0042778, 0.1085900, -0.1382730, -0.4584370, -0.4198630, -0.0939413, 0.0326470, 0.0024699, 0.0000841, 0.0024894, 0.0099668, 0.0552872, 0.0407054, 0.0802578, 0.1391490, 0.2404740, 0.1184250, 0.0847465, 0.2254810, -0.1394100, -0.2533980, -0.1248050, 0.2801330, 0.3943640, 0.2555240, -0.0439271, -0.2707520, -0.1110900, 0.0693892, 0.0595251, -0.0374515, -0.3819750, -0.2679430, -0.0047459, 0.0082537, 0.0185994, 0.0006032, 0.0017955, 0.0257635, 0.0633297, 0.0721785, 0.0653277, 0.2325690, 0.0494794, -0.0879069, 0.0507646, 0.1764400, -0.1694390, -0.4480990, -0.0909390, 0.2724170, 0.2703540, 0.2998000, -0.0307290, -0.1200420, -0.0303500, 0.1085210, 0.0328435, 0.0234083, -0.2135500, -0.2745000, -0.0938593, -0.0276777, 0.0067756, 0.0000315, 0.0039274, 0.0238924, 0.0543089, 0.1336510, 0.1091990, 0.1016470, 0.0018991, -0.0859369, -0.0314824, -0.1603490, -0.1548660, -0.3843870, -0.0783563, 0.2821850, 0.4416670, 0.1855050, 0.1681320, 0.1745680, 0.0737731, 0.3867920, 0.1163170, 0.0535695, -0.2739070, -0.4153930, -0.1721660, -0.0202936, 0.0043782, 0.0002595, 0.0048615, 0.0206716, 0.0274652, 0.2108620, 0.2800980, 0.0530207, -0.2386950, -0.2443200, -0.2159820, -0.2083830, -0.2050130, -0.4949630, -0.2755920, 0.2618700, 0.3716620, 0.4107750, 0.2134550, 0.2016870, 0.0928495, 0.2557700, 0.1559360, 0.0377127, -0.0527285, -0.2322730, -0.1354310, -0.0449155, 0.0104236, 0.0001433, 0.0046936, 0.0131997, 0.0407405, 0.1550420, -0.0655103, 0.0144815, -0.1246570, -0.1136060, -0.1246410, -0.1807180, -0.1863000, -0.2028750, -0.1476240, 0.2723110, 0.2316490, 0.5269310, 0.3345260, 0.1177510, 0.2283410, 0.0757105, 0.0618223, 0.0722044, -0.0684501, -0.2262920, -0.0876525, -0.0286889, -0.0005749, -0.0018886, 0.0065728, 0.0091438, 0.0342340, 0.0288225, -0.2171560, -0.2506840, -0.2440250, -0.0517099, -0.1590950, -0.2406600, -0.0396324, -0.0187803, 0.1500450, 0.0658068, 0.2762720, 0.3010530, 0.1398080, 0.0581938, -0.1595890, -0.2142040, -0.1922950, -0.0814267, -0.1088140, -0.2572740, -0.0601681, -0.0145795, 0.0001313, -0.0006573, 0.0066943, 0.0020271, 0.0148679, 0.0143475, -0.2054150, -0.3472990, -0.3460470, -0.0611124, -0.3015740, -0.2845250, -0.1034780, -0.0753593, 0.2918230, 0.3533470, 0.2855210, 0.1664690, 0.0814437, -0.0398900, -0.0545470, -0.1279030, -0.1531150, 0.0598156, -0.1177860, -0.1376400, -0.0889011, -0.0479861, -0.0069351, 0.0010745, 0.0025452, 0.0100846, 0.0070593, 0.0864763, -0.2069100, -0.3523820, -0.2782340, -0.1160370, -0.0635312, -0.0968885, -0.0132772, -0.1471430, 0.2233340, 0.2120080, -0.0327193, 0.0607507, -0.0007116, -0.1519940, -0.0909458, -0.0373992, -0.0121400, 0.0457927, -0.1244730, -0.0765694, -0.1367160, -0.0572958, -0.0123927, 0.0003798, 0.0013269, 0.0098963, 0.0477789, 0.0099184, -0.2184690, -0.5437270, -0.4078780, -0.1162130, -0.2548450, -0.2480240, -0.0702198, 0.1560270, 0.2074140, -0.0064841, -0.1474940, -0.0371912, -0.0433655, -0.1269280, 0.0642436, 0.0404720, 0.1130720, -0.0116894, -0.0974128, -0.0108626, -0.1062230, -0.0130622, -0.0093052, 0.0036239, 0.0009131, 0.0161136, 0.0500404, -0.0248985, -0.0275616, -0.2326650, -0.4039120, -0.3135280, -0.4246680, -0.1344030, 0.1091160, 0.0547317, 0.0895991, -0.0170672, 0.0981705, -0.0736729, 0.1232060, 0.0841474, 0.1224730, 0.0320002, 0.0621952, -0.0059545, -0.2682360, -0.0865467, -0.0795933, 0.0057936, -0.0035036, -0.0002637, 0.0086104, -0.0243364, -0.0277528, -0.0281026, -0.0543143, -0.0917227, -0.0718779, -0.2207950, -0.2701720, -0.2024330, -0.1218080, 0.0574714, 0.0770523, 0.1554480, 0.1348760, 0.0783983, 0.0899995, 0.1256420, 0.1946310, 0.0311048, -0.0894661, -0.2267830, -0.2754490, -0.0437454, -0.0428026, -0.0075821, 0.0000135, -0.0000224, 0.0031641, -0.0378956, -0.0127831, -0.0487531, -0.1198830, -0.0495082, 0.1023830, -0.0652667, -0.2855450, -0.2185810, -0.1753350, -0.0268879, 0.1008370, 0.2758190, 0.0374710, -0.0736464, -0.0525819, 0.0812720, 0.0801328, -0.0781416, -0.1239920, -0.2293100, -0.2539350, -0.0268244, -0.0245410, -0.0065234, -0.0002318, -0.0000997, -0.0005366, -0.0274980, -0.0153869, -0.0672440, -0.0812889, 0.0103589, -0.0120725, -0.0916965, -0.2608040, -0.1197160, -0.1408940, -0.0043434, 0.0322384, 0.0661240, -0.2111970, 0.0277123, 0.0988809, 0.1198070, -0.0377667, -0.1963870, -0.2117200, -0.2117810, -0.2328080, -0.1275460, -0.0194912, -0.0049928, -0.0000114, 0.0002396, -0.0000106, -0.0131995, -0.0303763, 0.0217603, 0.0438744, 0.0487508, 0.0703301, 0.0423163, -0.0257243, -0.0425592, -0.1675410, -0.1808050, 0.0283761, 0.1401370, -0.0283256, -0.0497949, -0.0368288, -0.0575277, -0.0862260, -0.0915638, -0.1744470, -0.0962007, -0.0796183, -0.0937661, -0.0241389, -0.0036242, 0.0000532, 0.0005439, -0.0002341, 0.0013179, 0.0158324, 0.0062817, 0.0427478, -0.0402110, -0.1191600, -0.1538990, -0.0239619, -0.0858728, 0.0005791, 0.0773348, 0.1259780, -0.0961705, -0.0075990, -0.1514350, 0.0336921, 0.1128030, -0.0021583, 0.0772616, -0.0849980, 0.0145198, 0.0416155, -0.0138342, -0.0143215, -0.0040688, 0.0002871, 0.0003243, 0.0004840, 0.0021802, 0.0286761, 0.1090180, 0.2122200, 0.2066620, 0.0084439, -0.0376041, -0.0721973, -0.0240862, -0.2003770, -0.2714390, -0.1197230, -0.0207895, 0.0697110, 0.1731690, 0.1523280, -0.0219316, 0.1502440, 0.1504660, -0.0028621, 0.0295500, 0.0621603, -0.0184167, -0.0107090, -0.0038086, 0.0001834, 0.0000721, 0.0006084, 0.0002745, 0.0002549, 0.0656441, 0.1657350, 0.1404590, 0.0920843, 0.2549390, 0.1937510, -0.0169056, -0.1170430, 0.0435120, -0.0047727, 0.1657990, -0.0285605, 0.0556013, 0.1691570, 0.0274557, 0.1111360, 0.0349185, -0.0529701, -0.1031070, -0.0693319, -0.0262075, -0.0037166, -0.0027394, -0.0001831, 0.0004366, 0.0000980, -0.0004073, 0.0006138, 0.0040524, 0.0506663, 0.0981769, 0.1393140, 0.1477040, 0.1669790, 0.1380330, 0.1005440, 0.0569803, 0.1174790, 0.1774760, 0.0867053, 0.1505860, 0.2315750, 0.2143230, 0.0655830, 0.1016420, 0.0840444, 0.0366571, 0.0044574, 0.0000521, -0.0002877, -0.0001454, 0.0001284, 0.0001074, -0.0004019, 0.0002746, 0.0001079, -0.0001577, -0.0001185, 0.0039740, 0.0268967, 0.0264637, 0.0060697, 0.0070723, 0.0093142, 0.0126161, 0.0203951, 0.0367404, 0.0344874, 0.0218716, 0.0276811, 0.0541549, 0.0213098, 0.0248371, 0.0320606, 0.0189296, 0.0010034, -0.0002572, -0.0001189, 0.0004224, 0.0004045, 0.0007118, 0.0004719, -0.0004212, -0.0001319, 0.0000985, 0.0003561, -0.0002506, 0.0000232, -0.0004226, 0.0003943, -0.0000767, 0.0001067, -0.0005138, 0.0004789, -0.0002999, 0.0001155, 0.0002093, -0.0000986, 0.0000289, -0.0002595, 0.0006632, 0.0003478, 0.0000353, 0.0003326, 0.0002336, -0.0003947, -0.0001647, -0.0006256, 0.0000639, 0.0009373, 0.0004530, -0.0005869, -0.0004452, 0.0005121, 0.0007868, -0.0000223, -0.0009134, -0.0013724, -0.0002846, 0.0000838, -0.0003479, -0.0006609, 0.0100918, 0.0188525, -0.0048678, -0.0006318, 0.0001417, 0.0001043, -0.0005717, 0.0002044, 0.0008156, 0.0013136, -0.0001883, 0.0004548, -0.0009178, -0.0000603, -0.0000060, 0.0006028, 0.0001580, -0.0000626, 0.0001408, 0.0003819, 0.0020838, 0.0020523, -0.0047169, -0.0071611, -0.0010060, 0.0113508, 0.0106259, 0.0301163, 0.0083135, 0.0423305, 0.0652867, 0.0554868, 0.0099045, 0.0083572, -0.0156929, -0.0119626, -0.0047635, -0.0038934, -0.0000612, -0.0000673, -0.0001770, -0.0002249, 0.0002933, 0.0004775, 0.0002009, 0.0001351, 0.0005343, -0.0352613, -0.0358684, -0.0539447, -0.0594823, -0.0324378, -0.0053723, -0.0135795, 0.0200866, 0.0893448, 0.1295460, 0.1529330, 0.1593020, 0.0374346, -0.0712062, 0.0210957, -0.0638950, -0.0671524, -0.0272488, -0.0336945, -0.0038459, -0.0056990, -0.0006627, -0.0002026, 0.0000371, 0.0001126, -0.0008433, -0.0013867, -0.0016070, -0.0412814, -0.0403987, -0.0257024, 0.0250655, 0.0050851, -0.0410929, -0.0434836, -0.0572193, 0.1149200, 0.1065450, 0.1632090, 0.1338580, 0.0488591, -0.0007872, 0.0506204, 0.0040902, -0.1392170, -0.0736136, -0.0783271, -0.1224330, -0.0373501, -0.0068926, 0.0000276, -0.0005200, 0.0000852, 0.0001878, -0.0002515, -0.0041143, -0.0294090, -0.0308947, 0.0115595, -0.0003042, -0.0354554, -0.0242048, 0.0025282, -0.0745094, -0.0591301, 0.1581370, 0.0743231, -0.0800148, -0.1691240, -0.1460390, 0.0091948, -0.0470282, 0.0787987, -0.0416069, -0.0420624, -0.1073440, -0.0792767, -0.0054296, -0.0019920, -0.0006308, -0.0001618, -0.0039469, -0.0024967, -0.0185161, -0.0805770, -0.0579123, 0.0479672, -0.0440466, -0.0384990, 0.0379910, 0.0101522, -0.0167400, -0.0864847, 0.1583250, 0.0907227, 0.0346633, 0.0241830, 0.0989714, 0.1534210, 0.0882362, 0.1590270, 0.0279735, -0.0252822, -0.0841784, -0.0864808, -0.0024140, -0.0056923, -0.0004304, 0.0004962, -0.0103253, -0.0240272, -0.0436629, -0.0631126, -0.0322670, -0.0400069, -0.1077590, 0.0601275, 0.2194580, 0.1789460, 0.0492716, 0.1545380, 0.0532619, 0.1359490, 0.2188690, 0.0229406, -0.0219155, 0.2649650, 0.0585567, 0.0460952, 0.0338234, -0.0552848, -0.1562020, -0.0708966, 0.0369346, -0.0020122, 0.0002647, 0.0010006, -0.0120782, -0.0212975, -0.0404470, -0.0863174, -0.0029045, 0.0345439, 0.0428295, 0.0846281, 0.0307846, -0.0153922, -0.0219279, -0.4016720, -0.0370998, 0.1802780, 0.1167470, 0.2141430, 0.0964341, 0.2048640, 0.0816543, 0.0258125, 0.0919443, -0.1179170, -0.1965090, -0.0803401, -0.0169444, -0.0031935, 0.0002278, 0.0008891, -0.0030578, -0.0036152, -0.0315101, -0.0533785, 0.0252075, 0.1069530, -0.0683067, 0.1278770, 0.0783788, 0.0908834, -0.0851546, -0.3704750, -0.2095250, 0.0479242, 0.0622858, -0.0286722, -0.0517203, 0.0555384, -0.0137369, 0.0985360, 0.1375820, -0.0409181, -0.1230600, -0.1006350, -0.0662283, 0.0020262, 0.0003649, -0.0002458, -0.0030047, 0.0052006, -0.0231297, -0.0443482, 0.0024734, 0.0317201, -0.0359248, 0.1331420, 0.1083640, -0.0379350, -0.2477330, -0.4526000, -0.3337790, 0.1114970, 0.0880233, 0.0444713, -0.2899380, -0.1701860, -0.1195310, 0.0619213, 0.0146756, 0.0433705, -0.1253310, -0.0634389, -0.0356953, 0.0011129, -0.0000830, 0.0007066, -0.0038784, -0.0074801, -0.0153200, 0.0096261, 0.0764199, -0.0222596, -0.0382493, 0.2039390, 0.1442190, -0.0511540, -0.3799450, -0.3692110, -0.1564330, 0.3034490, 0.0216390, -0.1069250, -0.2086960, -0.1809780, -0.0366574, -0.0508806, -0.0689148, 0.0588973, -0.0426463, -0.0470131, -0.0184033, 0.0004836, -0.0001180, 0.0001653, -0.0001855, 0.0144726, -0.0118211, -0.0239956, 0.1592960, 0.0355945, 0.1003290, 0.3355420, -0.1083790, -0.3282690, -0.4537090, -0.3331790, -0.0260704, 0.2543940, 0.1570830, -0.0768718, -0.2723460, -0.3631780, -0.0470605, -0.0653966, -0.0202297, 0.1820280, 0.0637236, -0.0191784, -0.0092688, 0.0005118, 0.0005126, -0.0000971, 0.0009313, 0.0151392, 0.0276264, 0.0248363, 0.1101060, 0.0559533, 0.1004220, -0.0732340, -0.2705010, -0.5144570, -0.4030410, -0.0108657, -0.0301462, -0.0491487, -0.0037179, -0.1716680, -0.3659880, -0.2607030, -0.1875170, 0.1144310, -0.0157250, 0.1071990, 0.1015650, 0.0418798, -0.0011635, 0.0004145, 0.0004566, -0.0007783, 0.0002145, 0.0114243, 0.0503640, 0.1029140, 0.0307193, 0.0240157, 0.0249664, -0.1139860, -0.4162130, -0.2063560, 0.0111662, -0.1711580, -0.1122670, 0.1146600, -0.0565703, -0.1698030, -0.3408620, -0.2677930, -0.1348710, 0.0002362, 0.0096523, 0.0531333, 0.1402940, 0.0107925, 0.0046330, 0.0002050, 0.0002839, 0.0002060, 0.0010155, 0.0059821, -0.0365240, 0.0090356, -0.1317370, -0.0809207, 0.1685140, -0.0445061, -0.2367430, -0.1191380, -0.1624810, -0.0808984, -0.0102216, 0.1073690, -0.0223306, -0.3721540, -0.4972430, -0.3060230, -0.0396950, 0.0066557, -0.1151820, -0.0322281, 0.0024950, -0.0195927, 0.0025696, 0.0002772, 0.0009674, 0.0004084, -0.0008851, -0.0172880, -0.0051069, 0.0077317, -0.1196500, -0.0173725, -0.0345923, -0.0610634, -0.1872350, -0.0984210, -0.1980710, 0.2476390, 0.1216260, 0.1564370, -0.2137990, -0.7365700, -0.6443210, -0.2425480, 0.0547020, -0.0338044, -0.1477520, -0.1135240, -0.0519701, -0.0022724, 0.0113650, 0.0018207, 0.0001459, 0.0004287, -0.0020248, -0.0319485, -0.0507458, -0.0463042, -0.0805663, 0.0349361, -0.0703719, -0.0860245, 0.0282445, -0.0911159, -0.0073165, 0.0348662, -0.0430422, -0.2520870, -0.6049600, -0.7817550, -0.4963390, -0.1374100, -0.0160499, -0.1094210, -0.0063752, -0.0982622, -0.0882737, 0.0499012, 0.0087782, 0.0000680, 0.0005418, -0.0005961, -0.0026117, -0.0392961, -0.1414010, -0.1537690, -0.1962650, 0.0086349, 0.0264164, 0.1997790, 0.1777370, -0.0302400, 0.0460157, -0.0604239, -0.1985280, -0.5076240, -0.6855720, -0.2814880, 0.0017408, 0.0838684, 0.1850050, 0.0832518, 0.0628969, -0.0308039, -0.0925749, 0.0547185, 0.0110682, -0.0005548, 0.0004596, -0.0002388, -0.0053602, -0.0396270, -0.1193990, -0.2479860, -0.0196252, 0.1257950, 0.1202890, 0.3085880, 0.2072580, 0.3400470, 0.2027010, 0.0363373, -0.2934990, -0.4631800, -0.0772899, 0.2459890, 0.2084450, -0.0029924, 0.2381120, 0.2003360, 0.1424200, -0.0302170, 0.0000288, 0.0619163, 0.0138926, -0.0003953, 0.0005733, -0.0001502, -0.0034430, 0.0039429, -0.0593930, -0.0857068, 0.0169716, -0.0463499, 0.0670503, 0.0884199, 0.1745680, 0.3004480, 0.3034600, 0.0666987, -0.0784153, -0.1036160, 0.1628990, 0.2457550, 0.0701827, 0.0146833, 0.0641193, 0.1796850, 0.1458190, 0.0859691, 0.0845270, 0.0568730, 0.0151144, -0.0000118, 0.0006848, -0.0013303, 0.0064119, 0.0503133, 0.0425712, 0.2136040, 0.0981856, 0.1777420, 0.1149140, 0.1425080, 0.3290300, 0.2271120, 0.2954650, 0.0895774, 0.0362849, -0.0255723, -0.0060351, 0.0420779, -0.0102477, 0.0648758, 0.1185540, 0.1119040, 0.1104710, 0.1738220, 0.0969669, 0.0341317, 0.0059050, -0.0003382, -0.0001786, -0.0002445, 0.0058625, 0.0136178, 0.0386462, 0.2924610, 0.1558950, 0.0241677, 0.2157140, 0.1731690, 0.0162514, -0.0234119, -0.0144081, -0.0012938, 0.1084180, -0.1485200, -0.1861620, -0.0907683, 0.1645670, 0.1708720, 0.0963151, 0.1290780, 0.1050760, 0.0821273, -0.0052315, 0.0044249, 0.0016557, -0.0007007, 0.0000392, -0.0008050, -0.0101971, -0.0512579, -0.0804960, 0.1299410, 0.1896380, 0.0555337, -0.0167197, 0.0996901, 0.0154985, 0.0684400, 0.1311550, 0.1201280, -0.0204674, -0.0653862, -0.0522512, 0.0144967, 0.0737484, 0.0999190, -0.0061798, -0.0165175, 0.0241984, 0.0048537, -0.0166247, 0.0067529, 0.0084602, 0.0006087, 0.0003263, 0.0004547, -0.0181851, -0.0372610, -0.0160030, 0.0972418, 0.0657901, 0.0233979, 0.0476790, 0.0322365, -0.0333429, -0.0022438, 0.0390029, -0.0548580, -0.0677616, -0.0864168, -0.2149750, -0.0250743, 0.0309606, -0.0517653, -0.1387890, -0.0703866, 0.0151225, 0.0079093, 0.0110517, 0.0078201, 0.0007564, -0.0001159, -0.0001248, 0.0001622, -0.0028034, 0.0049633, 0.0351167, 0.0567129, 0.0071975, 0.0305601, 0.0887524, 0.1084030, -0.0041930, 0.0029066, -0.0623658, -0.0962258, -0.1114880, -0.1803940, -0.1374240, -0.1214050, -0.1220450, -0.1250370, -0.0957869, -0.0613700, -0.0127379, -0.0013648, -0.0000327, 0.0007982, 0.0008579, -0.0002871, -0.0000354, 0.0000972, 0.0000514, 0.0001186, 0.0012829, 0.0115996, 0.0173718, 0.0042968, -0.0116426, -0.0250474, -0.0199702, -0.0090502, -0.0057853, -0.0272995, -0.0362076, -0.0326237, -0.0357506, -0.0425186, -0.0148159, 0.0054821, -0.0087655, -0.0245832, -0.0088625, -0.0004969, 0.0000398, -0.0007323, 0.0013686, -0.0000976, 0.0005873, -0.0002549, -0.0003114, -0.0002373, -0.0003162, -0.0000555, 0.0003838, -0.0002558, -0.0002222, -0.0001688, 0.0012593, 0.0001225, -0.0000907, -0.0006544, -0.0008893, -0.0006329, -0.0008662, -0.0020314, -0.0076864, 0.0005974, 0.0008942, -0.0009113, -0.0114699, -0.0026166, -0.0003033, 0.0006868, 0.0003326, -0.0000081, 0.0004600, 0.0002627, -0.0003899, 0.0000474, 0.0001640, 0.0002211, 0.0003370, 0.0004810, 0.0002232, 0.0000841, -0.0002889, -0.0006819, 0.0008611, 0.0015306, 0.0000215, -0.0000356, 0.0004341, -0.0001510, 0.0001680, 0.0000717, 0.0004513, -0.0000402, -0.0003739, 0.0002124, 0.0003203, -0.0000261, 0.0001986, 0.0005924, -0.0004544, 0.0001527, -0.0002237, 0.0003916, -0.0003492, -0.0001927, 0.0084582, 0.0154071, 0.0176889, 0.0088727, 0.0219222, 0.0220122, 0.0335608, 0.0466254, 0.0234616, 0.0237218, 0.0258269, 0.0207315, 0.0157583, 0.0083343, 0.0082675, 0.0066771, 0.0113866, 0.0073870, 0.0001607, 0.0000861, 0.0000438, 0.0002076, -0.0001248, -0.0001520, 0.0005117, 0.0002749, 0.0000920, 0.0007448, 0.0147128, 0.0392091, 0.0527918, 0.0349720, 0.0578890, 0.1101730, 0.1171200, 0.1275160, 0.1536050, 0.1459630, 0.1057650, 0.0954579, 0.0772920, 0.0029455, -0.0074101, -0.0085598, 0.0044711, 0.0062613, 0.0000688, 0.0004832, 0.0001952, 0.0004378, -0.0003753, 0.0004625, 0.0004128, 0.0029279, 0.0062710, -0.0147876, 0.0317963, 0.0289231, 0.0743466, 0.2809390, 0.2115850, 0.0484157, -0.0086292, 0.1483110, 0.1135260, 0.1711520, -0.0600159, -0.0965141, -0.0553015, -0.0463877, -0.0688123, 0.0038955, -0.0145311, -0.0016768, 0.0275642, 0.0001640, -0.0007197, -0.0001162, -0.0004498, 0.0003012, -0.0006744, -0.0004183, 0.0073282, -0.0674161, -0.0580495, -0.0593425, -0.0087383, 0.1219140, 0.0408594, -0.0584299, -0.1016000, -0.1038280, 0.1014030, 0.1745410, 0.0734575, -0.0898184, -0.0478836, 0.0757333, 0.0050190, 0.1001800, 0.0983538, 0.0505374, 0.0672569, 0.0130471, -0.0014816, 0.0000133, 0.0003179, 0.0001156, -0.0003236, -0.0048683, 0.0088659, -0.0370867, 0.0130901, -0.0449217, 0.0787026, 0.1143990, 0.0734530, 0.0522648, 0.0752942, 0.1871380, 0.0601360, 0.0710833, 0.1632890, 0.4324410, 0.1916390, 0.1365370, -0.0538773, -0.0673402, -0.0519922, -0.0810457, -0.0025900, -0.0345218, 0.0001949, 0.0002221, -0.0001636, -0.0002101, -0.0030745, -0.0020139, -0.0107204, -0.0211128, -0.0233385, -0.1769680, 0.1108580, -0.0677410, -0.1631940, -0.0503924, 0.0220477, 0.0915129, 0.2001080, 0.2143310, 0.3710620, 0.1494550, 0.1271830, 0.0456716, -0.2060260, -0.3006980, -0.2882970, -0.2334920, -0.1884510, -0.0268334, 0.0008135, 0.0008642, 0.0001178, 0.0014692, -0.0023963, -0.0746147, -0.0762955, -0.0459310, -0.0554713, -0.0070387, 0.0007607, -0.0076324, 0.0093260, -0.2078090, -0.2200230, -0.2782210, -0.2243910, -0.2967570, -0.2000690, -0.5636810, -0.7092970, -0.7831470, -0.8120340, -0.5800650, -0.4791740, -0.3755150, -0.2174680, -0.0890212, -0.0146445, 0.0025030, -0.0003912, 0.0161334, 0.0126278, -0.0305358, 0.0167763, 0.1282790, 0.1374000, -0.0367677, -0.0501374, -0.0358824, 0.0753691, 0.0859541, -0.3384200, -0.4831910, -0.7479100, -0.8857030, -1.0632700, -0.9632870, -0.8297240, -0.7737890, -0.6055520, -0.4860750, -0.3702370, -0.2953310, -0.1861440, -0.1158870, -0.0349302, 0.0038019, 0.0005077, 0.0250276, 0.0480014, 0.0436401, 0.2060680, 0.0564586, -0.0440639, -0.0571015, -0.0115958, -0.1428560, -0.0964588, -0.0323767, 0.0540614, -0.3680000, -0.2885490, -0.3787680, -0.5117850, -0.3476160, -0.3335350, -0.2875980, -0.2639160, -0.2845860, -0.1273360, -0.0613616, -0.0199324, -0.0017630, 0.0758863, 0.0929558, 0.0006327, 0.0199868, 0.0368920, -0.0228009, 0.1096130, -0.0724054, -0.0440571, -0.0296583, 0.0899872, -0.0522078, -0.2020790, 0.0428752, 0.1563420, 0.0454525, -0.1244030, -0.0101429, 0.1890500, 0.2314550, 0.0455778, 0.1643470, 0.2909850, 0.1122720, 0.1179390, 0.1606370, 0.1657260, 0.1537120, 0.0667759, 0.0195665, 0.0000591, 0.0117160, 0.1174010, 0.0392963, 0.0835475, 0.0499954, -0.0270717, -0.0758084, -0.0897780, 0.1679770, -0.0750296, 0.1290490, 0.0549011, 0.2509340, 0.2121690, -0.0601110, 0.4176720, 0.3107420, 0.4326380, 0.3702400, 0.2164810, 0.3450440, 0.3108200, 0.1910060, 0.1823020, 0.0843057, -0.0020054, 0.0033441, 0.0000626, 0.0032702, 0.0754506, 0.0853602, 0.0429269, 0.0254771, -0.0312458, 0.0317022, 0.1924910, -0.0036659, -0.1442100, 0.0747908, -0.1730530, -0.1485370, 0.1547270, 0.0954482, 0.0746065, -0.0089813, 0.1922850, 0.1086780, 0.0917595, 0.1194310, 0.2030520, 0.1689460, 0.0685223, 0.0975795, 0.0792698, 0.0135032, -0.0002223, 0.0016631, 0.0386991, 0.0327015, 0.0754435, 0.0908790, -0.0700846, 0.0585534, 0.1177830, -0.0142123, -0.0037006, 0.0891722, -0.1129850, -0.0648268, 0.0054486, 0.0190247, 0.0294819, -0.0743174, -0.0308897, 0.0203954, 0.1165860, 0.0413353, 0.0975278, 0.2993070, 0.1980270, 0.0803667, 0.0278199, -0.0058565, 0.0002367, 0.0002035, 0.0207914, 0.0394158, 0.0297002, -0.0915323, -0.2197060, -0.0975361, 0.0282230, -0.0365581, -0.0442545, 0.2089080, 0.0559951, -0.1427850, -0.0298655, 0.1614860, 0.0247179, -0.0629527, 0.0372828, -0.0894946, 0.1370910, 0.1214060, 0.1551200, 0.1293310, 0.0480848, 0.0147481, -0.0036535, -0.0000676, -0.0000345, -0.0012463, -0.0005783, 0.0262302, 0.0052451, -0.1619370, -0.0012545, -0.0749895, -0.0153770, -0.0934770, -0.0147623, 0.0790529, -0.1465020, -0.2306440, 0.0632444, 0.0374281, -0.1539640, -0.0390642, 0.0868689, 0.0725964, 0.2203300, 0.1404930, 0.0165252, 0.0060241, -0.0144747, 0.0397825, -0.0345587, -0.0021424, 0.0000734, -0.0005811, -0.0038916, 0.0226414, 0.0440579, -0.0715919, 0.0777277, -0.0226087, -0.0860472, -0.0428057, -0.0106667, -0.0034005, -0.1415930, -0.0807424, -0.0263846, -0.0135969, -0.0963523, 0.0450268, 0.0007098, 0.1185170, 0.0973385, 0.1260790, 0.0801857, 0.0001499, -0.0245328, 0.0524876, -0.0237195, -0.0054892, 0.0006442, -0.0002677, -0.0069503, 0.0093150, -0.0401159, -0.1022820, 0.0734479, -0.0439559, -0.0382471, -0.1467090, -0.1117880, 0.0550163, -0.0731029, -0.0463063, -0.0649454, -0.1353580, -0.1733670, -0.0145440, 0.0619050, -0.0655660, 0.0456094, 0.0028308, -0.0777240, 0.0165940, -0.0068715, -0.0049294, -0.0185370, -0.0140182, 0.0005087, 0.0002046, -0.0097107, -0.0256362, -0.0465496, 0.0122656, -0.1042720, -0.0564007, -0.0969364, -0.1633060, -0.0405814, -0.1248880, -0.0287360, 0.0057549, -0.0215104, -0.0608034, -0.0708625, 0.1395730, 0.0172024, -0.1914690, -0.1473180, 0.0649668, -0.1166360, -0.0048968, 0.0835519, 0.0130809, -0.0004809, -0.0007470, 0.0003888, 0.0158614, 0.0600374, 0.0614301, -0.0407400, -0.1597660, -0.0700306, -0.1189060, -0.1358420, -0.1069460, -0.0593483, 0.0883466, -0.0466604, 0.0999174, 0.0240241, 0.0395326, 0.0726065, 0.1616210, -0.1201140, -0.0049744, 0.0000312, -0.0554558, -0.1675730, 0.0255692, 0.1215100, 0.0341827, -0.0042602, -0.0005233, -0.0002420, 0.0001924, 0.0539451, 0.0724249, -0.0129018, -0.1439290, -0.0719281, -0.1721190, 0.0065413, 0.1549270, -0.0144708, -0.0868736, -0.0685138, -0.0415608, 0.0534368, 0.0597420, -0.0473018, 0.0160918, -0.0725700, -0.1019590, -0.1663420, -0.1755490, -0.1047840, 0.0632393, 0.0883500, 0.0574665, 0.0002313, -0.0000239, 0.0003221, 0.0002023, -0.0073830, -0.0180134, -0.0295281, 0.0075246, -0.0169965, 0.0722781, 0.0652524, 0.0146855, 0.0977906, 0.0783983, 0.0658587, 0.0226618, -0.0524602, 0.0741860, 0.0158751, 0.0949141, 0.0955863, -0.1307010, 0.0373501, -0.0190211, -0.0411685, 0.0678038, 0.0959043, 0.0827001, 0.0028461, 0.0002152, 0.0001501, -0.0001498, -0.0039146, -0.0156483, -0.0513492, -0.0529092, -0.1765480, -0.0206421, -0.0772547, 0.0313162, 0.0517129, 0.0462216, -0.1738270, -0.1671420, -0.3212090, -0.0865528, -0.0549346, 0.0228587, -0.1078660, -0.0636612, -0.0204684, -0.1335260, -0.0760680, -0.0275057, 0.0535549, 0.0402740, 0.0154995, 0.0001272, -0.0000831, 0.0004265, -0.0010490, -0.0083361, -0.0026107, 0.0230874, -0.0075996, -0.0046563, 0.0408414, 0.0191652, 0.0585511, -0.0064752, -0.0923073, -0.0317811, 0.1229040, -0.0190674, -0.0059925, -0.0650407, -0.1339370, 0.0312296, 0.0687996, -0.0544879, -0.0285128, 0.0118448, -0.0040156, 0.0333894, 0.0094591, -0.0006410, -0.0005056, -0.0005538, 0.0116024, 0.0132911, 0.0553973, 0.0993804, 0.0910254, 0.0605672, 0.0584867, 0.0598685, 0.1431560, -0.1087680, -0.0318754, -0.0960466, -0.2448020, -0.1401380, -0.0982595, -0.0164285, -0.1484320, 0.0356219, -0.0379625, -0.0736692, -0.0077108, 0.0534377, 0.0225033, -0.0014125, -0.0007641, 0.0002722, -0.0001380, 0.0001718, 0.0004352, 0.0008245, 0.0277569, 0.0072068, -0.0253778, -0.0360672, -0.0829428, -0.1179640, -0.0974979, -0.0351163, 0.0374707, -0.0323529, 0.0337812, -0.0576998, 0.0949625, 0.0311090, -0.0151682, 0.1004470, 0.0349932, 0.0434969, 0.0685043, 0.0602879, 0.0308896, -0.0004996, -0.0003593, 0.0003128, 0.0002619, -0.0000294, 0.0001556, -0.0003521, -0.0003281, -0.0002457, -0.0033762, -0.0053563, -0.0172128, -0.0102653, 0.0144540, 0.0369585, 0.0546696, 0.0362856, 0.0106328, -0.0007952, 0.0517872, 0.0069018, -0.0096919, 0.0753462, 0.0567830, -0.0018044, 0.0179169, -0.0015185, -0.0002514, -0.0002771, 0.0003427, -0.0002847, -0.0000742, 0.0005321, 0.0000414, 0.0002131, 0.0002780, -0.0001402, -0.0006744, -0.0046722, -0.0031635, 0.0038983, 0.0240762, 0.0083958, 0.0117402, 0.0088251, -0.0014342, -0.0110778, 0.0232602, 0.0010578, -0.0086820, 0.0194473, 0.0158937, 0.0034290, 0.0271945, 0.0071084, -0.0000365, 0.0002515, 0.0001507, 0.0002171, -0.0001542, -0.0004811, -0.0001070, 0.0000833, 0.0004043, 0.0010485, 0.0002332, -0.0004088, -0.0005490, -0.0005143, 0.0005226, 0.0004502, -0.0001189, -0.0003335, -0.0008941, 0.0001207, 0.0003815, 0.0004347, 0.0005649, -0.0007884, 0.0001237, 0.0004340, -0.0000637, 0.0002773, -0.0002437, 0.0003108, -0.0006576, 0.0005518, -0.0001155, -0.0000602, -0.0002288, -0.0002006, -0.0002056, -0.0002113, 0.0002472, -0.0008187, -0.0007305, -0.0003325, -0.0007460, 0.0000747, -0.0052837, -0.0057567, 0.0105082, -0.0006293, -0.0307772, -0.0182680, -0.0088175, -0.0064034, -0.0086109, -0.0052777, -0.0018960, -0.0003091, -0.0005799, -0.0002039, 0.0002809, 0.0000306, -0.0000413, 0.0000781, 0.0001194, 0.0001113, -0.0005956, 0.0005697, 0.0027170, -0.0002592, 0.0011224, 0.0209278, 0.0338724, 0.0192627, 0.0173997, 0.0371905, 0.0290192, 0.0381896, -0.0125250, -0.0142679, -0.0292734, 0.0141467, 0.0154090, 0.0072503, -0.0027558, -0.0012686, 0.0009769, 0.0000838, -0.0003256, -0.0000260, -0.0005722, 0.0003649, -0.0005340, -0.0013090, -0.0097802, -0.0036198, 0.0033019, 0.0154726, 0.0071867, 0.0427949, -0.0534812, -0.0748303, -0.0776046, -0.0536335, 0.0085952, -0.0080097, -0.0435904, -0.0832141, -0.1695030, -0.1347730, -0.1206210, -0.0190659, -0.0040644, -0.0085285, -0.0084661, 0.0008747, -0.0002370, -0.0001526, -0.0006383, -0.0003564, 0.0004853, -0.0015625, 0.0015204, 0.0452599, 0.1095100, 0.1022410, 0.0948413, 0.0658345, -0.1033380, -0.1147440, -0.0672480, 0.0093041, -0.0663951, -0.1514450, -0.0786148, -0.0330710, -0.0220275, -0.0804128, -0.0525705, -0.1145780, -0.0279035, -0.0187547, -0.0462420, 0.0026206, -0.0026547, 0.0003420, -0.0004007, 0.0002554, 0.0005882, -0.0066470, 0.0206033, 0.1001210, 0.1051930, 0.0360256, 0.1904120, 0.1336150, 0.0367708, -0.0763787, 0.0149525, 0.0951322, -0.0378153, -0.0400950, -0.1064720, -0.1250410, -0.0166497, -0.0529902, -0.0929474, -0.0851325, -0.0972271, -0.0735948, -0.0771160, -0.0165081, -0.0160068, -0.0000818, -0.0003849, -0.0000508, 0.0003353, -0.0012411, -0.0098096, -0.0398618, -0.0873631, -0.0726192, 0.0739865, 0.0059741, -0.0217388, -0.0104957, -0.0709870, -0.1848670, -0.0986993, -0.1423380, -0.1052710, 0.0494660, -0.0630954, -0.1693970, -0.1828820, -0.1830910, -0.2751220, -0.1559720, -0.2007630, -0.0908945, -0.0293784, -0.0017402, 0.0000031, -0.0042624, 0.0067475, -0.0343533, -0.0091810, -0.0409766, 0.1169900, 0.1358250, -0.0561808, -0.0365366, -0.1252980, -0.1387210, -0.0509389, -0.1229260, -0.1192030, -0.1405100, -0.0531193, -0.1159380, -0.2354030, -0.1329330, 0.0219254, 0.0351177, -0.1218470, -0.2404490, -0.0924054, -0.0570577, -0.0240374, -0.0022764, -0.0044753, -0.0003484, 0.0222011, 0.0227187, 0.0683975, 0.0992685, 0.0725561, 0.0172705, -0.0440768, -0.0104844, 0.0351727, 0.0421099, -0.1846560, -0.2939910, -0.1550890, -0.1618870, -0.1304230, -0.1413230, -0.0002726, -0.0488774, -0.0145889, -0.0171770, -0.2779570, -0.1416700, -0.0560760, -0.1019530, -0.0373624, -0.0092329, 0.0001291, -0.0010801, 0.0336963, 0.0580088, 0.0408534, 0.0349742, -0.0251692, -0.1198340, -0.0691173, 0.0939786, 0.0980271, -0.0265478, -0.2073370, -0.3300840, -0.2122190, -0.0879962, -0.1662260, 0.0308992, -0.0501924, 0.0432058, -0.0015139, 0.0863255, -0.1934300, -0.1505480, -0.0940206, -0.1235400, -0.0409060, -0.0021621, 0.0000762, 0.0004970, 0.0074255, -0.0350423, -0.0042487, 0.0904806, 0.1014190, 0.1597210, -0.0957311, 0.0628287, -0.0408957, 0.0667621, -0.0980571, -0.3082050, -0.2471970, -0.2689660, -0.0958672, 0.0770230, 0.1384040, 0.1552520, -0.0826061, 0.0395306, -0.0803464, -0.1061510, -0.1541480, -0.0775226, -0.0248938, -0.0009183, 0.0001906, -0.0017336, -0.0088223, -0.0920748, -0.0714148, 0.1116630, 0.2149970, 0.1533950, -0.0580420, -0.0189691, -0.0366700, 0.0057858, 0.0407719, -0.1748690, -0.3261970, -0.2079420, -0.0261282, 0.1342310, 0.0518022, 0.1108630, 0.0955245, 0.1230810, 0.0376522, -0.1145220, -0.2043130, -0.1019370, -0.0270513, -0.0004568, 0.0000307, 0.0008099, 0.0044813, -0.0377384, 0.0227070, 0.2182350, 0.0990974, -0.0423475, 0.0394589, -0.0732483, -0.0533298, 0.0527400, -0.0070571, -0.2866560, -0.4715650, -0.2764050, 0.0362394, 0.1653390, 0.1186930, 0.2351190, 0.1609840, 0.1550450, 0.0795252, -0.0910171, -0.0792745, -0.0667901, -0.0229041, 0.0007601, -0.0008937, -0.0016816, 0.0035496, -0.0905187, 0.0649103, 0.1610330, 0.0140211, 0.0501062, 0.0837770, 0.0721623, 0.1851430, 0.1908340, -0.1054400, -0.4878700, -0.4417140, -0.0927540, 0.1120360, 0.3054780, 0.0912419, -0.0126596, 0.1357390, 0.1717210, 0.1711510, 0.0187217, -0.0322969, -0.0116630, -0.0041017, 0.0050986, -0.0008624, -0.0040192, -0.0028693, -0.0629998, 0.0837567, 0.0847960, 0.0246664, 0.0650819, 0.1234390, 0.0588689, 0.1401770, 0.1056690, -0.2161640, -0.3740360, -0.1891920, 0.0643471, 0.3763520, 0.2496580, 0.2500210, 0.1557650, 0.2827840, 0.1319660, 0.2293640, 0.0391491, -0.0960139, 0.0186213, 0.0118915, 0.0005913, 0.0000406, -0.0072487, -0.0072987, 0.0384805, -0.0059022, -0.1318950, 0.0100909, -0.0030527, 0.0773907, 0.1123890, 0.1228030, 0.1162660, -0.3800250, -0.4982030, -0.2182280, 0.3472750, 0.3102420, 0.2503700, 0.1402170, 0.3085170, 0.2776730, 0.1200210, 0.1327980, -0.0737801, -0.1015650, 0.0216943, 0.0558286, 0.0018809, 0.0003814, -0.0038298, -0.0251419, -0.0131107, -0.0032651, -0.0530242, 0.0684820, -0.0018113, -0.0728873, 0.0392069, 0.0391695, 0.0262391, -0.4594810, -0.5952050, 0.1011000, 0.6972610, 0.4679020, 0.2041660, 0.1964150, 0.2322010, 0.2073820, 0.1541320, 0.0033252, -0.0826816, -0.0439283, 0.0458935, 0.0477968, 0.0046684, -0.0004419, -0.0012776, -0.0241783, -0.0794765, -0.0536376, -0.0276501, 0.0258081, -0.1592130, 0.0709808, 0.0058289, 0.0154048, -0.2582960, -0.6274540, -0.2965790, 0.3622350, 0.7648340, 0.3414340, 0.1165230, 0.3077930, -0.0798372, 0.0816844, 0.1790930, -0.0463774, -0.0822049, 0.0120086, 0.0987941, 0.0227803, -0.0007743, -0.0004045, -0.0005238, -0.0196910, -0.1066030, -0.0800374, -0.0692757, -0.0019007, 0.0658029, -0.0013996, -0.1089650, -0.2183680, -0.2976140, -0.3776990, -0.1481620, 0.3874650, 0.4985640, 0.2559620, 0.3188700, 0.2054980, 0.0369481, 0.0397556, 0.1151510, -0.1069560, -0.0199534, 0.0721871, 0.0804549, 0.0039482, 0.0022165, 0.0000982, -0.0006925, -0.0223535, -0.0706661, -0.0559492, -0.0178684, 0.1024320, 0.1059680, -0.0859252, -0.1437610, -0.1762260, -0.1867600, -0.2927100, -0.0300900, 0.3886410, 0.5259760, 0.4658810, 0.0772325, -0.0463133, 0.0199635, -0.1659910, -0.0154198, -0.1212940, 0.0528601, 0.0882812, 0.0378636, 0.0156403, 0.0004338, -0.0000159, -0.0017101, 0.0023979, -0.0405297, -0.0827520, 0.0060028, -0.0159617, 0.0183589, -0.1085320, -0.4140230, -0.3763740, -0.2765100, -0.0525160, -0.0541773, 0.0875505, 0.0503212, 0.3008640, 0.1787830, 0.0888534, -0.0023413, -0.1594300, -0.0973386, -0.1433250, -0.0118009, 0.1421580, -0.0000647, 0.0067072, 0.0000697, -0.0000054, -0.0005131, 0.0365664, 0.0005066, -0.0431054, 0.0121800, -0.1299140, -0.2856600, -0.0589979, -0.1687230, -0.1289120, -0.1354550, -0.1331320, 0.1183230, -0.0057832, 0.0349372, 0.2606810, 0.2299150, 0.0726943, 0.0563873, -0.0622446, -0.0891325, -0.1400930, 0.0089173, 0.1241070, -0.0384860, -0.0044998, -0.0002042, -0.0003899, -0.0000579, 0.0166190, -0.0074178, -0.0509059, -0.1169650, -0.1378440, -0.2581790, -0.0018233, -0.0747188, -0.1019480, -0.1150110, -0.0847414, -0.1190490, -0.0379645, 0.0463037, 0.1275210, 0.0825135, -0.0352338, -0.0168735, -0.0267923, -0.0374741, -0.0547004, -0.0342335, 0.0591923, -0.0090802, -0.0175468, 0.0001999, -0.0001374, -0.0003991, -0.0285672, -0.0583385, -0.0891753, -0.1634770, -0.1879200, -0.1156310, -0.1138980, 0.0451036, 0.0345070, -0.0674988, -0.0002664, -0.1118530, -0.0361683, -0.1343140, -0.1932400, -0.1058620, -0.0315266, 0.0697607, 0.0397558, 0.0426284, -0.0253287, -0.0374820, 0.0250351, -0.0146877, -0.0105418, 0.0003076, -0.0000526, -0.0000100, -0.0292231, -0.0572806, -0.0732620, -0.1062620, -0.0950347, -0.1302250, -0.1033440, 0.0517926, -0.0410549, -0.0879881, -0.1436000, -0.0000908, -0.0245108, -0.0767127, -0.0024990, 0.0468365, 0.1048050, 0.1946390, 0.0880222, 0.0866171, -0.0240046, -0.0539518, -0.0058685, 0.0150388, 0.0017664, 0.0004381, 0.0004460, -0.0001028, -0.0046463, -0.0030454, -0.0186412, -0.0157602, 0.0194494, -0.0312058, -0.0131564, -0.0364400, -0.1862990, -0.0451507, 0.0408787, -0.0032066, 0.2168790, 0.1786220, 0.0723650, 0.0449334, 0.1547730, 0.0305709, 0.1397500, 0.0746948, -0.0322269, -0.0485416, -0.0280094, 0.0014794, 0.0020300, -0.0004013, 0.0004004, 0.0006215, -0.0000239, -0.0005490, 0.0040939, 0.0244787, 0.0466766, 0.0547590, 0.0791500, 0.1217860, 0.0137905, -0.0240115, 0.0092457, 0.0493862, 0.0923617, 0.0583818, 0.0288897, 0.0321245, 0.0857986, 0.0464063, 0.0687320, 0.0797585, 0.0325261, 0.0017714, 0.0003754, -0.0005666, -0.0001503, 0.0004553, 0.0000316, -0.0004331, -0.0001765, 0.0009322, -0.0002415, -0.0006242, 0.0003161, 0.0033952, 0.0038737, 0.0041580, 0.0125637, 0.0085257, 0.0052226, 0.0203799, 0.0216404, 0.0207780, 0.0133084, 0.0171782, 0.0353438, 0.0364687, 0.0297817, 0.0472032, 0.0354264, 0.0031933, -0.0004585, 0.0005186, 0.0000650, -0.0004961, -0.0004861, 0.0001073, 0.0003780, -0.0003606, 0.0001421, -0.0001219, 0.0005121, 0.0003375, 0.0003548, -0.0002628, 0.0005614, -0.0000072, -0.0011250, -0.0021914, -0.0002236, -0.0001321, 0.0000256, -0.0003820, -0.0002008, 0.0001814, -0.0003974, -0.0005236, -0.0004505, -0.0002989, 0.0000657, 0.0000417, 0.0002412, -0.0000967, 0.0007212, 0.0005640, 0.0003691, -0.0001738, -0.0001334, -0.0001674, -0.0056208, -0.0092093, -0.0133442, -0.0036531, -0.0029240, -0.0019368, -0.0050070, -0.0088890, 0.0013842, 0.0039074, -0.0019025, -0.0057931, -0.0044979, -0.0037390, -0.0015285, -0.0007990, -0.0054209, -0.0059080, 0.0000444, 0.0002176, 0.0002488, -0.0004294, 0.0000468, 0.0004901, 0.0001660, -0.0002300, -0.0000261, -0.0012009, -0.0094458, -0.0229457, -0.0236732, -0.0157108, -0.0283649, -0.0458853, -0.0682146, -0.0872381, -0.0850674, -0.0726085, -0.0582049, -0.0105464, 0.0284520, -0.0077793, 0.0013057, -0.0007249, -0.0061227, -0.0071571, -0.0015373, -0.0012077, -0.0004207, -0.0000830, 0.0001265, 0.0005720, 0.0004128, 0.0001716, -0.0005074, -0.0035830, -0.0330049, -0.0406724, -0.0386434, -0.1130800, -0.1076700, -0.0925590, -0.0712518, -0.0538797, -0.1210330, -0.1151160, -0.2028020, -0.1115090, 0.0005691, -0.0331398, -0.0219836, 0.0277470, 0.0607517, -0.0104195, -0.0275108, -0.0012978, -0.0011988, 0.0002382, -0.0003955, 0.0005419, 0.0017367, 0.0021601, 0.0065795, -0.0133266, -0.0512602, -0.0465135, -0.1127990, -0.1840780, -0.0744890, 0.0123536, -0.1000400, -0.1608490, -0.0033170, 0.1410790, 0.0773084, 0.0857010, 0.0855802, -0.0484443, -0.0366688, 0.0223057, 0.0980906, 0.0798657, 0.0321671, 0.0406775, 0.0173136, -0.0011221, -0.0002904, -0.0001894, 0.0005357, 0.0011826, -0.0028396, -0.0557945, -0.0397978, -0.0382383, -0.2208940, -0.2121390, -0.1499410, 0.0061404, -0.0080975, -0.1864310, -0.1394640, -0.1180180, -0.0272693, 0.0588209, -0.0794869, 0.1034970, 0.0989582, -0.0379717, 0.0250868, 0.0193018, 0.0024700, 0.0401789, 0.0032220, -0.0020382, -0.0006155, 0.0003033, 0.0130186, -0.0464804, -0.0387982, 0.0136870, 0.1090260, 0.0705335, -0.0387022, 0.0249771, 0.0781374, 0.0665938, -0.0193181, -0.0911619, -0.1517960, -0.1990480, -0.0628493, 0.0114670, 0.0427384, -0.1114940, -0.0168165, -0.1037660, -0.0579459, 0.0528468, 0.0462690, 0.0630476, 0.0125507, -0.0044047, -0.0004846, -0.0033855, 0.0042354, -0.0481678, -0.0563650, 0.0356926, 0.1302710, -0.0451472, 0.2044450, 0.0271651, 0.0567089, 0.0482239, -0.0488681, -0.0581309, -0.1682010, -0.1558670, -0.0558552, 0.0508391, 0.1208390, 0.0318172, -0.0241064, -0.0589076, -0.1152970, -0.0814355, 0.0207032, 0.0939866, 0.0340704, -0.0011606, 0.0000794, -0.0148489, -0.0083971, 0.0333927, -0.0217640, -0.0051180, -0.0442011, -0.0959389, -0.0474283, -0.1716850, -0.1962410, -0.1743690, -0.0207740, -0.2243780, -0.2942690, -0.1938690, 0.0800883, 0.0438412, 0.0422889, -0.0235629, -0.1215010, 0.0338815, -0.0196438, -0.0992766, 0.0734523, 0.1006470, 0.0449300, 0.0099702, 0.0000665, -0.0155055, 0.0170689, 0.0586718, -0.1425270, -0.1370230, -0.0429840, 0.0981467, -0.0295329, 0.1112310, 0.0943960, 0.0545254, 0.0144383, 0.0033806, -0.1161540, -0.0087505, 0.1541430, 0.0421976, -0.0567259, -0.1141590, 0.0416619, -0.0222107, 0.0804187, 0.0555434, 0.0641430, 0.0639113, 0.0086028, -0.0913351, -0.0006585, -0.0152132, -0.0389754, 0.0876753, -0.0190220, -0.0561658, -0.0610211, -0.0523409, 0.0219760, 0.0369916, 0.1340720, 0.0622525, 0.0634680, -0.3534600, -0.4512540, -0.1158180, -0.1723680, -0.0127235, -0.0077218, -0.1318000, -0.0566554, -0.0403173, 0.1766010, 0.2619540, 0.1207200, 0.0674409, -0.0091241, -0.0213945, -0.0001405, -0.0149478, -0.1057860, -0.1118850, 0.0015269, -0.0047245, 0.0370094, -0.0624258, 0.0562314, 0.0402724, -0.1290010, -0.1386150, -0.2456140, -0.4730650, -0.5435510, -0.2463700, 0.0062356, -0.0063474, -0.0909708, 0.0614781, 0.0535990, 0.0552756, 0.2580970, 0.2029850, 0.1520900, 0.1102430, 0.0322285, -0.0034917, 0.0004719, -0.0032942, -0.0730264, -0.1614750, 0.0605242, 0.1357590, 0.2811750, 0.0738987, -0.2190120, -0.1707440, 0.0555160, -0.1888810, -0.0026851, -0.0244393, -0.1464650, -0.2024290, -0.2198360, -0.2632540, 0.0644546, 0.1257910, 0.2059750, 0.1557800, 0.1174400, 0.1305750, -0.0529305, -0.0238685, -0.0230278, -0.0229640, 0.0006241, -0.0021028, -0.0457387, -0.1174150, 0.0916722, 0.0941751, 0.1345980, 0.3080190, 0.0942422, 0.1376370, 0.1566180, 0.3192620, 0.3471070, 0.1992410, -0.0187666, -0.2241420, -0.3549260, -0.0821017, 0.1638960, 0.2139750, 0.0918484, -0.2152530, -0.1573980, -0.2211780, -0.2414900, -0.0826218, -0.0150287, -0.0020770, 0.0000115, 0.0024033, -0.0303290, -0.0197965, 0.1570950, 0.0994824, 0.1777950, 0.2726990, 0.4150010, 0.3001470, 0.4274820, 0.2273610, 0.3665980, 0.4893220, 0.1111040, 0.0240598, -0.0781097, 0.0961708, -0.1894950, -0.2285730, -0.1863330, -0.1910070, -0.3419400, -0.4072860, -0.2443410, -0.0804543, -0.0113354, -0.0004526, -0.0001391, 0.0090151, 0.0020901, 0.0103019, 0.0966892, 0.1653340, 0.1372430, 0.1132330, 0.3259420, 0.2528470, 0.2273340, 0.0320623, 0.4341810, 0.3470710, 0.2910490, 0.0366383, 0.2082870, -0.0198417, -0.1310100, -0.1973230, -0.3609250, -0.2818560, -0.2989810, -0.2007380, -0.1524670, -0.0619653, -0.0030427, -0.0007418, 0.0004059, 0.0045608, 0.0183115, -0.0089250, -0.0633423, -0.0738287, -0.1033950, 0.0600858, -0.0056035, 0.0083335, 0.0079693, 0.1741640, 0.3658900, 0.3221410, 0.1975290, 0.1352000, -0.0128034, -0.1999930, -0.0598488, -0.2020750, -0.2532350, -0.1530550, -0.1894480, -0.1939070, -0.0973178, -0.0461289, -0.0193220, -0.0013745, 0.0001433, 0.0012744, 0.0210390, -0.0466549, -0.1913250, -0.2399280, -0.1755110, 0.0143695, 0.0705451, 0.0243248, 0.0266147, 0.2421910, 0.3765420, 0.3409960, 0.2091500, 0.0330539, 0.1512510, -0.1144810, -0.2456340, -0.2680530, -0.2685240, -0.1142450, -0.1490960, -0.2118620, -0.1973850, -0.1211110, -0.0311600, -0.0013976, -0.0015826, -0.0008494, 0.0114587, -0.0493299, -0.2123600, -0.1789550, -0.1329400, -0.2638980, -0.2347650, -0.2587470, 0.1657300, 0.3621200, 0.2466390, 0.0932628, -0.0406011, 0.0411342, -0.0321369, -0.1755780, -0.2581980, -0.1145910, -0.0330977, 0.0520212, 0.0551234, -0.1026860, -0.1026550, -0.0603760, -0.0175426, -0.0017179, 0.0004934, -0.0035659, 0.0039935, -0.0287945, -0.0943066, 0.0323753, -0.1439270, -0.4538720, -0.6619090, -0.6166300, -0.4378140, -0.4495790, -0.4351040, -0.1609160, -0.0362132, 0.1149290, 0.0202567, -0.0485192, 0.2807300, 0.2087520, 0.0269659, 0.1426770, 0.1199940, 0.0503022, -0.0268081, -0.0147869, -0.0017851, -0.0001626, -0.0001351, 0.0005006, 0.0028999, -0.0006827, 0.0504227, 0.0931466, 0.0156462, -0.1307200, -0.3335020, -0.4490280, -0.6977700, -0.7269880, -0.7575830, -0.1931200, -0.0396393, 0.0386535, 0.1235170, 0.1251350, 0.2807910, 0.0831538, -0.0577849, 0.0256315, 0.1317920, 0.0953275, 0.0064035, 0.0176578, -0.0029869, 0.0002314, 0.0002815, 0.0000972, 0.0018813, 0.0159068, 0.1015900, 0.0666315, 0.1770830, 0.1766010, -0.0273085, -0.0756731, -0.1829100, -0.1253570, -0.2044670, -0.2786500, -0.1362670, 0.0718417, 0.1147990, 0.2357820, 0.2442260, -0.0950027, -0.0641720, 0.2090920, 0.1974730, 0.0542751, 0.0598340, 0.0341383, -0.0020785, 0.0001331, -0.0003729, 0.0004677, 0.0023789, 0.0107393, 0.0905765, 0.0397654, 0.1954720, 0.1345760, 0.1098280, 0.2140110, 0.1274150, 0.1524860, -0.0541012, 0.1824630, -0.0122424, -0.2150950, -0.1167320, 0.0867059, 0.1646140, -0.0545943, 0.0565415, 0.1160190, 0.1911340, 0.1010100, 0.0667470, 0.0499158, 0.0080998, -0.0004843, 0.0003110, -0.0002031, 0.0096476, 0.0325241, 0.0869744, 0.1060060, -0.0286909, 0.0424762, 0.3585030, 0.2175110, 0.2345690, 0.1593970, -0.0516082, 0.2070100, 0.1611970, -0.0222881, -0.1673640, -0.0133316, 0.0563978, -0.0027230, 0.1682270, 0.1735960, 0.1985450, 0.1403650, 0.0481533, 0.0316712, 0.0043804, 0.0002183, 0.0005741, 0.0005815, 0.0068229, 0.0294406, 0.0894795, 0.0416757, 0.0819820, 0.1295500, 0.2027170, 0.1719240, 0.3050390, 0.2383200, 0.1224210, 0.0852335, 0.1714290, -0.0592205, -0.0719375, 0.0231129, 0.1514320, 0.2338030, 0.3058430, 0.2705730, 0.1789000, 0.1238640, 0.0076411, -0.0056893, -0.0039370, 0.0000772, -0.0002709, -0.0001718, 0.0011058, -0.0195057, -0.0180654, 0.0384381, 0.0555350, 0.0727249, 0.0417920, 0.1064910, 0.1116140, -0.0170588, 0.0537269, 0.2266000, 0.0693340, 0.0316383, 0.1214210, 0.0768930, 0.0988409, 0.2921510, 0.2447520, 0.1481580, 0.0600006, 0.0527980, 0.0147290, -0.0032381, -0.0036112, 0.0001418, 0.0003758, -0.0000319, -0.0005848, -0.0001357, 0.0141667, 0.0674562, 0.1004830, 0.0325070, -0.0465342, -0.0896874, -0.0687029, 0.0601470, 0.1676880, -0.0433009, 0.0441217, 0.0795777, 0.1156120, 0.1380890, 0.0492488, -0.0573761, 0.0559966, 0.0434786, -0.0153580, 0.0070632, 0.0002487, 0.0004224, 0.0000593, -0.0003741, 0.0001279, 0.0005258, 0.0004957, -0.0001966, 0.0003849, -0.0008301, 0.0008747, 0.0094183, 0.0076153, 0.0011823, -0.0146238, 0.0144616, 0.0249649, -0.0155850, 0.0221232, 0.0083303, -0.0417520, -0.0223121, 0.0228027, 0.0027774, 0.0013828, -0.0433557, -0.0174771, -0.0026458, -0.0001743, 0.0004291, 0.0000316, 0.0001832, 0.0001584, 0.0009150, -0.0003807, 0.0005252, -0.0001825, 0.0005104, -0.0004580, 0.0005696, -0.0002925, -0.0002945, -0.0001320, -0.0002019, -0.0004631, -0.0000486, -0.0001951, -0.0005107, -0.0003508, -0.0002850, -0.0004241, 0.0000317, 0.0002299, -0.0004474, 0.0000498, -0.0005206, -0.0007725, 0.0000277, -0.0000361, -0.0004208, -0.0000871, -0.0001246, 0.0003277, -0.0001161, -0.0002524, 0.0001947, 0.0000273, 0.0002257, -0.0000966, 0.0000969, 0.0007139, 0.0002169, -0.0002025, 0.0004687, -0.0292245, -0.0483831, -0.0035517, -0.0003443, 0.0000002, -0.0013724, -0.0014364, 0.0003776, -0.0001855, -0.0006363, 0.0002835, -0.0001212, -0.0003820, -0.0001570, -0.0002544, 0.0001753, -0.0004747, 0.0005089, 0.0009095, 0.0003356, 0.0002538, 0.0001180, 0.0134108, 0.0292387, 0.0130452, 0.0127743, 0.0147048, -0.1940120, -0.0829524, -0.1847650, -0.1821200, -0.1130660, -0.0672307, -0.1100310, -0.0172841, 0.0087057, 0.0049002, 0.0014279, 0.0006532, 0.0003245, -0.0006069, -0.0002156, 0.0000934, 0.0006637, -0.0001819, -0.0001253, 0.0003507, 0.0102187, 0.0129837, 0.0227525, 0.0496012, 0.0821367, 0.1307580, 0.2554280, 0.1383110, -0.0772143, -0.0385399, -0.0938300, -0.2211270, -0.1924630, -0.1426180, -0.1223060, -0.0148376, 0.0023862, 0.0272870, 0.0200833, 0.0050958, 0.0007395, -0.0000628, 0.0003464, 0.0000299, -0.0006517, -0.0012880, -0.0002620, -0.0063823, -0.0540722, -0.0131787, 0.0271719, -0.0165972, -0.0057692, 0.1149430, 0.1752500, 0.0929389, -0.2788690, -0.1753810, -0.1920150, -0.0576531, 0.0530222, 0.0044197, -0.1099720, -0.0047934, -0.0169202, 0.0253994, 0.0154110, 0.0336927, 0.0121033, 0.0005163, 0.0000347, 0.0000703, -0.0001443, 0.0001781, 0.0038783, 0.0194954, -0.1215010, -0.0983694, 0.0087393, 0.0623732, 0.0609571, 0.0231522, 0.0292287, 0.0062777, -0.0486621, -0.1735610, -0.2962180, 0.1784580, 0.1570380, 0.0291763, 0.0029786, -0.1156010, -0.0711404, -0.0250938, -0.0300576, 0.0271448, 0.0231763, -0.0002536, -0.0002848, 0.0002586, 0.0007422, 0.0094590, 0.0488539, 0.0678326, 0.0080181, 0.0151309, 0.0783241, 0.1197030, 0.2490490, 0.0245956, 0.0079546, 0.0009949, -0.2905410, -0.1210400, -0.0145190, 0.1253250, 0.0228393, -0.1302030, -0.0133486, -0.0374970, -0.1076420, -0.0599686, -0.0315787, -0.0006314, 0.0090756, 0.0010113, -0.0002663, -0.0000803, 0.0002763, 0.0386868, 0.0484215, 0.1104390, 0.1474400, 0.1166500, 0.0697975, 0.1594540, 0.0345531, -0.1292190, 0.0157495, -0.0989872, -0.0746829, -0.1677850, 0.0422120, 0.0246180, 0.1318280, 0.0338005, 0.1553870, -0.0177254, -0.0551791, 0.0052475, 0.0190288, -0.0036878, 0.0115063, -0.0021146, -0.0009337, 0.0003615, -0.0004133, 0.0309062, 0.0200376, 0.1324760, 0.1584040, 0.1789120, 0.1132340, 0.0496644, 0.0393313, -0.0178074, 0.0548036, -0.1397820, -0.0306022, -0.0730587, 0.1477290, 0.2814540, 0.2433000, 0.1614850, 0.2436600, 0.0675175, 0.0470272, 0.0519431, 0.0502702, -0.0110155, -0.0011388, -0.0018857, -0.0001985, 0.0003729, 0.0008299, 0.0188127, 0.0015937, 0.0577397, 0.1804880, 0.1611370, 0.0289039, -0.0440593, 0.0221913, -0.0467057, -0.2002220, -0.1002180, -0.1613540, -0.2234170, -0.0347617, 0.3257490, 0.2376160, 0.2870140, 0.2140940, 0.0945889, 0.1408600, 0.1163500, 0.0489849, -0.0004588, -0.0059705, 0.0013237, -0.0000870, 0.0010291, 0.0000897, 0.0095599, 0.0076497, 0.0472381, 0.1559310, 0.1401790, 0.0958662, 0.0209145, 0.0153754, 0.0118247, -0.1300420, -0.0941935, -0.2802990, -0.1852790, 0.0085257, 0.1695780, -0.0443860, 0.2731910, 0.1298050, 0.1825150, 0.1408340, 0.1249990, 0.0426976, 0.0081156, -0.0023703, 0.0039727, -0.0000028, 0.0000185, -0.0001489, -0.0006538, 0.0205154, 0.0498594, 0.0865441, 0.1125150, 0.1243400, 0.2812270, 0.1054480, -0.0911077, 0.0219466, 0.1280960, -0.1290000, 0.0080532, 0.1896900, -0.0111277, -0.0705544, 0.1300770, 0.1798470, 0.1595910, 0.1357670, 0.1078800, 0.0597527, 0.0290117, 0.0105245, 0.0047891, -0.0027259, 0.0005393, -0.0000986, 0.0001852, 0.0149326, 0.0382002, 0.0500910, -0.0139034, 0.0324004, 0.0767922, -0.0067209, -0.0177493, -0.1613310, 0.0220699, -0.0296016, 0.0550861, 0.0734553, 0.2192650, 0.1204460, 0.0410155, 0.1974430, 0.1749390, 0.1535150, 0.0905062, 0.0586653, 0.0319439, 0.0060692, -0.0018620, -0.0036974, 0.0000350, 0.0000041, 0.0001238, 0.0058178, 0.0212171, 0.0336661, -0.0477944, 0.0432302, 0.0469148, 0.0623364, 0.2568580, 0.1466990, 0.1204270, 0.3308580, 0.1804700, 0.0031426, 0.1024350, 0.0608163, 0.2847350, 0.1912980, 0.1406640, 0.1143920, 0.0999922, 0.0677655, 0.0269950, 0.0064964, 0.0004137, -0.0001605, 0.0003507, 0.0009738, 0.0021159, 0.0003740, 0.0071650, 0.0034988, 0.0596377, 0.1722150, 0.0673984, 0.1246680, 0.2043440, 0.3129630, 0.0676409, 0.2397610, -0.0054511, -0.0162172, 0.0597230, 0.0929752, 0.2348730, 0.2553470, 0.1022390, 0.1371250, 0.0933378, 0.0899505, 0.0308924, 0.0049308, -0.0012269, 0.0000282, 0.0000418, 0.0042140, 0.0022341, 0.0019468, 0.0115158, 0.0569566, 0.0854109, 0.1517030, 0.0460811, 0.0409419, 0.2435560, 0.2461790, 0.0351678, -0.0056811, -0.1916180, 0.0378223, 0.0157736, 0.0377226, 0.1905910, 0.2280820, 0.1470870, 0.1497240, 0.0920627, 0.0956847, 0.0423825, -0.0003444, 0.0014476, 0.0006282, -0.0006322, 0.0013166, 0.0041116, 0.0137880, 0.0344611, 0.0884401, 0.1182730, 0.1292390, 0.0814255, 0.0915953, 0.2351070, 0.2619750, 0.1866060, 0.1764510, -0.2256950, -0.1001020, 0.0476760, 0.1535340, 0.1556030, 0.1959890, 0.1833380, 0.1480070, 0.1304830, 0.1278440, 0.0355355, 0.0078435, 0.0032620, 0.0015258, 0.0002356, 0.0005249, 0.0051192, 0.0118639, 0.0579990, 0.0875268, 0.0417006, 0.0198462, -0.0705731, 0.1045580, 0.1807450, 0.3281200, 0.1822830, 0.1135690, -0.3578390, -0.3569180, 0.0247895, 0.0382556, 0.1034610, 0.2134160, 0.1609410, 0.0658236, 0.0622402, 0.0650814, -0.0307587, 0.0428964, 0.0070744, 0.0007444, 0.0001228, 0.0004922, 0.0039831, 0.0123680, 0.0442893, 0.0247656, 0.0559653, 0.0321499, -0.0380258, 0.1255570, 0.3597330, 0.5250280, 0.3723090, 0.1929780, -0.4929170, -0.4479190, 0.0638306, -0.0290719, -0.0977467, 0.0660421, 0.0756735, -0.0672612, -0.0387196, -0.0676391, -0.1144870, 0.0009889, 0.0042594, 0.0006046, -0.0001558, 0.0006442, -0.0144117, 0.0033699, 0.0269842, 0.0398053, -0.0392671, -0.0335202, -0.0755588, -0.0632483, 0.2422570, 0.3077650, 0.2730040, 0.0152394, -0.4634980, -0.4916550, -0.3547510, 0.0395188, -0.0716003, -0.1557570, -0.0896083, -0.0250517, -0.0717829, -0.1379530, -0.0751860, -0.0160473, 0.0059353, 0.0001427, 0.0004270, 0.0000398, -0.0110153, -0.0176856, -0.0022084, 0.0887679, -0.0754634, 0.0437257, -0.0775413, -0.0913708, 0.2087460, 0.1947860, 0.1663250, -0.0424275, -0.3125780, -0.2221740, -0.2285260, -0.1549790, -0.4124580, -0.3775580, -0.0023052, -0.0241499, -0.0652858, -0.0917925, -0.0441984, -0.0107327, 0.0015365, -0.0002287, 0.0003587, 0.0001448, -0.0001359, -0.0390425, -0.0856236, -0.2143260, -0.3010080, -0.2637890, -0.3467490, -0.0984250, 0.0987780, 0.1873160, 0.0463403, -0.0747629, -0.1273580, -0.2588190, -0.2684780, -0.1450330, -0.3005500, -0.1446030, -0.1530540, -0.1239830, 0.0281995, 0.0270227, -0.0458380, -0.0483463, 0.0009538, 0.0003537, 0.0000135, -0.0002524, -0.0001360, -0.0183953, -0.1190890, -0.2547570, -0.2671790, -0.0901387, -0.1093510, -0.0093902, 0.2183890, 0.1692970, -0.0119750, 0.0544162, 0.0007903, -0.2188800, 0.0541017, -0.1275830, -0.1578390, -0.0279972, -0.0693599, 0.0153136, 0.0393669, 0.0596038, -0.0174297, -0.0206170, -0.0001617, 0.0002444, -0.0001045, 0.0004279, 0.0008625, 0.0087215, -0.0159788, -0.0239509, -0.0404593, 0.0649800, 0.1852220, 0.0931044, 0.1895670, 0.3153120, -0.0940844, -0.0548687, -0.1516270, -0.1183160, 0.2011170, 0.0357619, 0.0793993, 0.0171522, 0.0397153, 0.0619569, 0.0607160, 0.0611987, 0.0345115, 0.0064460, -0.0002346, 0.0000432, 0.0003166, -0.0005634, 0.0007599, 0.0077788, 0.0113466, 0.0159441, 0.0245887, 0.0585013, 0.1039820, 0.0735481, 0.0507754, 0.1994720, 0.2100910, 0.2170640, 0.2607690, 0.1523660, 0.1704270, -0.0738774, -0.0743892, 0.0441519, 0.0391235, 0.0674249, 0.0832189, 0.0256266, 0.0175626, 0.0022375, 0.0002128, 0.0004137, -0.0003182, 0.0003192, 0.0000446, 0.0000025, 0.0049577, 0.0097330, 0.0079782, 0.0020882, 0.0105534, 0.0084525, 0.0203661, 0.0496629, 0.1443110, 0.1464460, 0.0565375, 0.0553502, 0.0947873, 0.0807596, 0.0933604, 0.0576754, 0.0103825, 0.0039874, 0.0031549, 0.0000222, 0.0001111, 0.0000222, 0.0005206, -0.0000767, 0.0001159, 0.0000952, 0.0004229, 0.0005460, 0.0001517, -0.0002367, -0.0001304, 0.0009488, 0.0012169, 0.0017424, 0.0038012, 0.0076544, 0.0571837, 0.0679348, 0.0457593, 0.0116257, 0.0041810, 0.0164210, 0.0198778, 0.0073539, 0.0035160, 0.0010832, 0.0001234, -0.0000129, 0.0002558, -0.0001147, 0.0002312, -0.0001950, -0.0004667, 0.0004290, 0.0007682, 0.0003656, 0.0004652, -0.0003716, -0.0002086, -0.0004731, 0.0003652, -0.0001155, 0.0011825, 0.0015477, 0.0035136, 0.0044655, 0.0016958, -0.0000699, -0.0007660, -0.0000111, 0.0000980, -0.0005056, -0.0007138, 0.0002179, -0.0001189, -0.0004084, 0.0001223, 0.0002380, -0.0005143, 0.0000599, -0.0003398, -0.0002172, -0.0001971, 0.0002839, 0.0002465, -0.0001679, 0.0003879, 0.0000012, 0.0005663, 0.0003146, 0.0002841, -0.0000799, 0.0005602, 0.0003847, 0.0001944, -0.0003092, 0.0005729, -0.0009014, 0.0004263, 0.0004497, -0.0002376, -0.0002044, 0.0005505, -0.0000272, 0.0002353, 0.0001283, -0.0006959, -0.0001244, -0.0002963, 0.0003387, 0.0004245, -0.0006229, -0.0001243, 0.0001946, -0.0041989, -0.0064938, -0.0089837, -0.0052302, -0.0156998, -0.0033546, -0.0022917, -0.0039938, -0.0176930, -0.0407420, 0.0061303, 0.0017885, -0.0028070, -0.0031382, -0.0064080, -0.0033578, -0.0019458, -0.0016218, -0.0000023, -0.0000421, 0.0001764, 0.0006107, -0.0002169, 0.0003946, 0.0005082, 0.0000359, -0.0006286, 0.0002235, -0.0014042, -0.0105946, 0.0067634, 0.0585459, 0.0175887, 0.0073023, -0.0087526, -0.0362720, -0.0816218, -0.2029340, -0.1440810, -0.0337543, -0.0688949, -0.0876908, -0.0288244, -0.0139667, -0.0137716, -0.0029993, 0.0094473, 0.0065700, 0.0003508, -0.0004370, -0.0000446, -0.0003632, 0.0010378, 0.0001447, -0.0007994, 0.0033670, 0.0086786, 0.0233884, 0.0723481, 0.0981400, 0.1058750, 0.1536420, 0.1134950, -0.0056192, -0.1288700, -0.2211030, -0.2813170, -0.2361930, -0.1977180, -0.1641290, -0.1342370, -0.0542011, 0.0189383, 0.0087439, 0.0208348, 0.0116373, 0.0004137, -0.0000439, 0.0000941, -0.0001301, 0.0038599, 0.0003941, -0.0030876, 0.0522617, 0.1114640, 0.1217340, 0.0700634, 0.0752582, -0.0081108, -0.0172811, 0.0051109, 0.0293931, 0.1166460, -0.0539074, -0.1785250, -0.2281370, -0.0334903, -0.1515940, -0.1114780, -0.0372664, 0.0529919, 0.1189920, 0.0817218, 0.0220514, -0.0120275, -0.0114779, -0.0004304, -0.0004545, 0.0006748, 0.0014054, 0.0142482, 0.0016884, -0.0289016, 0.0614546, 0.0598622, 0.1079300, 0.1633300, 0.0471169, 0.0680210, 0.0734861, -0.0568178, -0.0258002, 0.0683967, -0.1564990, -0.0102975, -0.1049140, -0.1579640, 0.0659937, 0.0050063, 0.0642991, 0.0284704, -0.0281278, -0.0358140, -0.0142245, -0.0005574, -0.0004544, -0.0117969, 0.0584705, 0.1012350, 0.0663875, 0.0936680, -0.0187693, -0.0234077, 0.1812860, 0.1043220, -0.1569520, -0.0384274, -0.1389930, -0.0455979, -0.1886410, -0.0794747, -0.1183090, -0.1257190, -0.0523323, -0.2455820, 0.0949544, -0.0718734, -0.0740523, 0.0224122, 0.0473072, 0.0350974, -0.0004053, 0.0002679, 0.0032329, -0.0002162, 0.0749208, 0.1317810, 0.1583360, 0.0358099, 0.0105990, 0.0772740, 0.0479181, -0.1045240, -0.1266120, 0.0036440, 0.1164590, -0.0149880, -0.2249520, 0.0264138, -0.0714242, 0.0317060, 0.1821600, 0.0316830, 0.0992532, 0.0346820, -0.1791640, -0.0441081, 0.0254541, 0.0158300, -0.0000858, -0.0062626, 0.0015134, -0.0091636, -0.0198941, 0.2059540, 0.0623030, -0.1048400, -0.0992261, -0.0559250, -0.1380930, -0.0315633, -0.0823736, -0.0209292, -0.1285610, 0.1144080, -0.0302983, -0.1586540, -0.0206016, -0.0857321, -0.0187404, 0.0294509, -0.0670363, 0.0287939, 0.0320434, -0.1420280, -0.0766881, -0.0345939, -0.0006392, 0.0001966, 0.0036764, 0.0040392, -0.0128640, 0.1106570, 0.2372710, 0.0345696, 0.0043984, 0.0030223, 0.0833345, -0.0440179, 0.0213832, 0.3539980, 0.2007890, 0.3546990, 0.1877150, 0.0220519, 0.0586817, 0.0291390, -0.0594289, -0.1072080, -0.2111390, -0.0691217, 0.0096069, -0.1370810, -0.0941534, 0.0299089, 0.0494107, -0.0001741, 0.0000024, -0.0005811, -0.0446097, 0.0243957, 0.3728730, 0.3955140, 0.2809530, 0.2842470, 0.3395470, 0.3779220, 0.2837910, 0.2557850, 0.5183760, 0.1173930, 0.0467423, -0.0119905, 0.0093474, -0.0244775, -0.1025490, -0.2045020, -0.1236240, -0.1736510, -0.0665965, -0.0773322, 0.0232600, 0.0893893, 0.0144408, 0.0000080, 0.0009861, -0.0061797, -0.0306419, 0.0976203, 0.2835030, 0.2289950, 0.1709850, 0.2727940, 0.3260630, 0.1869050, 0.3262350, -0.0199412, -0.3505810, -0.2439650, -0.2438690, -0.2609190, -0.0665671, -0.0947799, -0.0046626, -0.0876496, -0.1655150, -0.1853060, -0.2535450, -0.1704290, -0.0296008, 0.0144205, 0.0009131, 0.0004545, 0.0019505, 0.0017439, -0.0179974, 0.0297108, 0.0064309, -0.1515230, 0.0271990, 0.3083790, 0.0672109, -0.1311600, -0.3883880, -0.5181350, -0.8852310, -0.5142160, -0.1721960, -0.0538566, 0.0497482, -0.0684315, 0.0322069, -0.0575032, -0.1313750, -0.2187550, -0.3379750, -0.0873728, 0.0936737, 0.0474106, 0.0126765, -0.0001730, 0.0012162, 0.0108105, -0.0720707, -0.1591620, -0.2519900, -0.3092870, -0.3286510, -0.2419510, -0.4517370, -0.5021090, -0.8026580, -0.7963690, -0.2143690, -0.0019966, -0.2403620, 0.0121685, -0.0439581, -0.0338533, -0.0948679, 0.0081052, -0.2957340, -0.1415390, -0.1040030, 0.0718753, 0.0945934, 0.1001790, 0.0185807, -0.0000275, 0.0012695, 0.0141697, -0.1122780, -0.3529160, -0.5906350, -0.6887080, -0.7952970, -1.0024200, -1.1201300, -0.8975850, -0.5592880, -0.2698610, -0.1691750, -0.3189560, -0.1549280, -0.0257979, -0.1672210, -0.0307567, 0.0517836, -0.0207518, 0.0272207, 0.0311304, 0.0517692, 0.0930764, 0.0513785, 0.0751185, 0.0018089, -0.0001099, -0.0003757, 0.0039707, -0.1053770, -0.4270180, -0.7527730, -0.7653910, -0.8972240, -0.9383990, -0.5347280, -0.1290330, 0.0564248, 0.0918949, 0.0421316, -0.0599562, -0.1376860, 0.0431077, -0.0644814, -0.1868950, -0.0668021, 0.0811233, 0.0257895, -0.0861665, -0.0478359, 0.0888096, 0.0464190, 0.0454159, 0.0114829, -0.0002492, 0.0002143, 0.0012391, -0.0432153, -0.3576270, -0.6046520, -0.4112970, -0.3413370, -0.2357030, 0.2140490, 0.3519740, 0.0309094, -0.0466705, 0.2298780, -0.0348086, -0.1354000, -0.0616504, -0.1440390, -0.0263718, 0.0373652, -0.0367219, 0.1436650, 0.0280089, -0.0214110, 0.0136021, 0.0842458, 0.0557914, 0.0202381, 0.0001187, -0.0000349, 0.0026000, -0.0280670, -0.1368100, -0.1369690, -0.1020180, -0.0759511, 0.1934500, 0.2191920, 0.2348860, -0.0078922, 0.1645480, 0.2395680, -0.1176540, -0.1354910, -0.0416404, 0.0351076, -0.0181328, -0.0256937, -0.1088400, 0.1445530, -0.0428357, -0.0509837, -0.0167051, 0.2121940, 0.0783115, 0.0191894, -0.0001823, -0.0008128, 0.0019116, -0.0238157, 0.0334034, 0.1046640, 0.1544340, 0.2604030, 0.1605340, 0.0333657, -0.0339162, -0.0106547, 0.1351340, -0.0398692, -0.0856528, 0.1146250, 0.0408533, 0.0046811, 0.0743026, 0.1007000, -0.0300047, 0.1424910, 0.1158380, 0.1856670, 0.2212110, 0.1404520, 0.0204856, 0.0099957, -0.0000126, -0.0006715, 0.0100437, -0.0017903, 0.1247390, 0.1761130, 0.1800490, 0.2184430, 0.2346090, 0.0301085, -0.0849371, 0.1940870, 0.1212660, 0.3291620, 0.1843190, 0.0458083, 0.0797526, 0.0131440, -0.1374650, 0.0588112, -0.1542070, -0.0954005, 0.0159830, 0.1462220, 0.1440100, 0.0964690, 0.0286016, 0.0016943, -0.0000094, -0.0003934, 0.0314850, 0.1166360, 0.1505640, 0.2045400, 0.1782030, 0.1525920, 0.0851518, 0.2400730, 0.0322627, 0.1121510, 0.0846033, 0.1273450, 0.0877965, 0.0970574, 0.0927981, -0.1607280, -0.0175391, -0.0246983, -0.0659834, -0.0954264, -0.0442900, 0.1163900, 0.0383185, 0.0252291, 0.0142270, -0.0003235, -0.0010040, -0.0000511, 0.0615793, 0.0457998, -0.0688246, 0.0932728, -0.0033426, -0.1703350, -0.0626219, 0.1608290, 0.0202147, 0.1261850, 0.0797589, 0.0113575, 0.1290030, 0.1952100, 0.1498150, 0.0633812, 0.1940320, 0.0502634, -0.1139950, -0.1129860, 0.1151670, 0.1966540, 0.1065510, 0.0531699, 0.0046634, -0.0001934, 0.0000956, 0.0004424, 0.0611441, 0.0464545, -0.0808198, 0.0056079, -0.0046837, 0.1386200, 0.0212464, 0.1254530, 0.0576588, 0.0740859, 0.0729478, 0.1973190, 0.1366280, 0.1445750, -0.1090000, -0.0327153, 0.1683570, 0.0802402, 0.0706712, 0.1225000, 0.1448830, 0.1390850, 0.0656715, 0.0330489, 0.0046941, -0.0000257, 0.0004522, 0.0003479, -0.0005256, 0.0297989, 0.0525407, 0.0776040, 0.0408373, 0.0083382, -0.0785028, 0.1440860, 0.0359915, 0.1322740, -0.0189073, -0.0017060, -0.0959548, 0.1104570, -0.0730269, 0.0131917, 0.0691275, 0.0189022, 0.0329033, 0.0929062, 0.0763111, 0.0614112, 0.0464087, 0.0313077, 0.0044632, -0.0001139, -0.0003374, -0.0000881, -0.0037918, -0.0038581, 0.0851795, 0.0334016, 0.0622986, 0.0036101, 0.0233894, 0.0781484, -0.0554728, -0.0738403, -0.0810067, 0.0370184, 0.0551714, 0.1145450, 0.0296933, 0.3155960, 0.2273430, 0.1612970, 0.0593910, 0.1162440, 0.0831673, -0.0040491, 0.0609653, 0.0230170, 0.0051353, 0.0006286, -0.0000171, -0.0000807, -0.0001725, 0.0040019, 0.0557838, 0.0120667, 0.0580765, 0.1227760, 0.1710300, 0.0860555, -0.0356445, 0.0054531, 0.1311300, 0.0885108, 0.1255830, 0.3445760, 0.2021860, 0.1267970, 0.1290630, 0.1200730, 0.0372718, -0.0136865, -0.0095859, -0.0274094, -0.0031547, 0.0050058, 0.0062441, 0.0002331, -0.0000471, -0.0002826, -0.0001016, -0.0006347, -0.0047290, -0.0823453, -0.0581998, 0.0054100, 0.0523545, 0.0295034, -0.0286154, -0.0884267, -0.0435344, 0.1084740, 0.1165590, 0.0879798, -0.1563080, -0.1704930, -0.0530109, 0.0745716, 0.0024536, -0.0463212, -0.0236747, -0.0029334, -0.0003995, 0.0000147, -0.0005002, 0.0006969, 0.0000841, 0.0004116, -0.0001956, 0.0002315, 0.0006593, 0.0008920, 0.0004886, -0.0022101, -0.0015315, 0.0077190, 0.0282239, 0.0033979, 0.0001507, 0.0234595, -0.0226424, -0.0424948, -0.0279319, -0.0114521, -0.0446177, 0.0017347, 0.0027650, -0.0073446, -0.0255585, 0.0002607, -0.0004108, 0.0004942, 0.0000674, -0.0006077, 0.0001915, -0.0000108, -0.0001462, 0.0001447, -0.0000102, 0.0001935, 0.0000213, -0.0000913, -0.0000933, -0.0002520, -0.0004569, -0.0000232, 0.0002438, -0.0011694, -0.0004781, 0.0002424, -0.0005603, 0.0000641, 0.0000917, 0.0000161, 0.0003682, -0.0001529, 0.0005657, 0.0000708, -0.0002916, 0.0000159, 0.0002097, -0.0006576, -0.0002875, 0.0004872, 0.0000972, -0.0001353, -0.0001907, -0.0003144, 0.0019607, 0.0018867, 0.0002667, -0.0022484, -0.0031325, 0.0010236, -0.0075955, -0.0068233, -0.0047905, -0.0069601, -0.0127702, -0.0091996, -0.0036410, -0.0034596, -0.0085588, -0.0107548, -0.0008709, 0.0014856, -0.0002720, 0.0002232, 0.0006347, -0.0002294, -0.0001059, -0.0002756, -0.0006207, -0.0002112, -0.0007052, 0.0003424, 0.0008970, 0.0004432, 0.0031466, 0.0175827, 0.0286248, 0.0173006, -0.0213277, 0.0139684, 0.0332380, 0.0338902, 0.0213554, 0.0262072, -0.0015626, -0.0087225, 0.0013494, -0.0085264, -0.0137304, -0.0003381, 0.0023248, 0.0007594, 0.0004496, 0.0000885, 0.0001565, 0.0000013, -0.0001388, -0.0003609, -0.0032961, -0.0254261, -0.0171228, -0.0231123, -0.0436086, -0.0127757, -0.0780139, -0.0820970, -0.1213260, -0.1395260, -0.0731147, 0.0137242, 0.1328080, 0.0773640, 0.0279034, -0.0094618, -0.1255460, -0.0210647, 0.0143926, 0.0014787, 0.0139614, -0.0050011, -0.0014991, 0.0002589, -0.0002295, -0.0001441, 0.0005033, -0.0027981, -0.0069936, -0.0175600, -0.0137912, -0.0049949, -0.0191456, -0.0612786, -0.0451943, -0.1034850, -0.0457362, 0.1120370, 0.1154720, -0.0348729, 0.0899541, 0.1641740, 0.1080990, 0.0049468, -0.0054818, -0.1464290, -0.0573704, -0.0656342, -0.0830768, -0.0330262, -0.0100528, -0.0014106, -0.0000900, -0.0002105, 0.0007499, -0.0165296, -0.0014227, -0.0120268, -0.0331721, -0.0935864, -0.1890180, -0.2760150, -0.1071920, -0.1868590, -0.2282380, -0.1179450, -0.0739004, 0.0072561, -0.0569983, -0.0556274, 0.2520100, 0.2861710, 0.0314257, -0.0448173, -0.1519910, -0.1324310, -0.0952063, -0.0546049, -0.0145692, -0.0017282, -0.0002557, 0.0004256, -0.0110358, -0.0077634, -0.0321939, -0.1620890, -0.1541470, -0.1758880, -0.3569060, -0.4204000, -0.2106980, -0.0859124, -0.2515820, -0.2477700, 0.0375988, -0.1211450, -0.0020357, 0.0306853, 0.1695780, 0.0871956, -0.0502059, -0.1815730, -0.2896910, -0.2616740, -0.2403740, -0.0645325, -0.0135310, 0.0002554, 0.0000271, -0.0048924, -0.0052808, -0.0411022, -0.1111230, -0.2863680, -0.2620150, -0.3042070, -0.3531020, -0.3099550, -0.3114840, 0.0554110, -0.0392496, 0.0014132, -0.0534569, -0.0136647, 0.2117250, 0.1042980, 0.0475443, 0.0074465, 0.1253460, 0.1431310, -0.0260896, -0.2459980, -0.1715550, -0.0630457, -0.0024220, -0.0010887, -0.0018513, -0.0025940, 0.0005536, -0.0472596, -0.1547060, -0.3463490, -0.3098800, -0.4242290, -0.3939710, -0.2481210, -0.1277660, 0.0519327, 0.0831125, 0.0877770, -0.1483320, -0.1616800, 0.1996100, 0.1746710, -0.1152100, 0.0228181, -0.0574054, -0.0681159, -0.1477340, -0.1024060, -0.1188580, -0.0880786, -0.0373677, -0.0019845, -0.0004608, -0.0054414, -0.0086129, -0.0378673, -0.1822520, -0.3706960, -0.3029390, -0.3390290, -0.3753550, -0.1138650, 0.0763802, 0.1649000, 0.1862270, 0.1942300, -0.0484956, 0.0118019, -0.0295371, -0.2803450, -0.2465830, -0.2776370, -0.2388440, -0.0994305, -0.1327300, -0.2187500, -0.2043870, -0.1740310, -0.0717821, -0.0375737, -0.0008810, -0.0010648, -0.0284327, -0.0572339, -0.0854204, -0.0930550, -0.0824164, -0.1966350, -0.2316980, -0.1880520, 0.0343507, 0.1410360, 0.2360290, 0.1146210, 0.1583250, 0.1194100, -0.1345580, -0.4572190, -0.4654400, -0.2549250, -0.3380370, -0.1601320, -0.2958220, -0.3242350, -0.2784770, -0.1472540, -0.0490274, -0.0136337, 0.0002863, -0.0035812, -0.0200024, -0.0925236, -0.0575743, -0.0998153, -0.0697508, -0.1189830, -0.1521600, -0.0619777, 0.1604210, 0.1162070, -0.0266771, 0.0047426, 0.0446829, 0.0172200, -0.1667860, -0.2877220, -0.2911720, -0.0206351, -0.0378733, -0.1952420, -0.2922510, -0.3603500, -0.2121070, -0.0032234, -0.0510218, -0.0049428, -0.0002633, -0.0025083, -0.0260859, -0.0621843, -0.0136495, -0.1336480, -0.1187510, -0.1375170, 0.0684050, 0.1930370, -0.0074957, -0.0019010, -0.0693876, -0.0416587, 0.2019420, -0.0401399, -0.0052545, -0.1336950, -0.0397826, 0.0590295, 0.0448226, -0.0672291, -0.2512740, -0.3799090, -0.1829420, 0.0525192, -0.0633600, -0.0048092, -0.0009874, -0.0030265, -0.0161846, -0.0020753, -0.0211570, -0.1356890, -0.0512915, 0.1054160, 0.1678090, -0.0330175, -0.0393777, -0.1206230, 0.0217849, 0.2692710, 0.2300300, -0.0077147, -0.0157548, 0.1514940, 0.0059397, 0.0118291, -0.0890832, -0.0887543, -0.2584250, -0.2605120, -0.0704425, 0.0507388, 0.0118255, 0.0146945, -0.0004886, -0.0047408, -0.0082817, 0.0781137, 0.1263540, -0.1163460, 0.0166878, 0.0937361, 0.0621949, 0.0512470, -0.0092320, -0.0114278, -0.1248640, 0.0414712, 0.0685501, -0.1438970, 0.0802534, -0.0074031, -0.0120250, -0.1464420, -0.1421320, -0.2493400, -0.1548500, -0.0815338, 0.0289809, 0.1608280, 0.0738605, 0.0014727, -0.0002436, -0.0058105, 0.0026679, 0.1207930, 0.1507470, 0.0049274, 0.0588730, -0.0121839, 0.1271290, 0.1856430, 0.1297430, 0.0166697, -0.0826405, 0.1916710, 0.0251013, -0.0053257, 0.2957890, 0.1028280, -0.2087310, -0.0209374, -0.2415380, -0.1450760, -0.1461290, -0.1151160, 0.0546572, 0.2286820, 0.0694193, 0.0216645, 0.0000650, -0.0025831, 0.0055534, 0.0895025, 0.1131340, 0.1429070, 0.1402120, 0.1717020, 0.0079864, 0.1042620, 0.1383680, 0.2403850, -0.0049655, 0.0248138, 0.1929020, 0.1894700, 0.3061960, 0.0857276, -0.1697190, -0.1411980, -0.1522090, 0.1470370, 0.1895400, 0.0436420, 0.1349720, 0.2915920, 0.1605680, 0.0414976, -0.0008338, -0.0004947, 0.0030364, 0.0608420, 0.0583834, 0.1262650, 0.0874014, 0.0146326, 0.0772668, 0.0632946, 0.2460090, 0.1284900, 0.2304680, 0.0303511, 0.2041180, 0.3274560, -0.0046055, -0.2158440, -0.1928690, -0.1740610, -0.0308921, 0.1477350, 0.1686570, -0.0190567, -0.0062290, 0.1729650, 0.0339164, -0.0006924, -0.0001996, 0.0000687, -0.0073259, 0.0364940, 0.1003650, 0.0909036, -0.0317813, -0.0071468, 0.2520250, 0.2788190, 0.2256230, -0.0318030, 0.1366110, 0.1400040, 0.2110250, 0.1102750, -0.1230120, -0.1654700, -0.1355540, -0.0189914, -0.0844311, 0.0209910, 0.1703760, 0.1019890, 0.1194350, 0.1304690, -0.0099001, 0.0100832, 0.0002760, -0.0106632, -0.0182277, -0.0660037, 0.0889896, 0.0401613, -0.1092940, -0.1586650, -0.1511790, -0.0394519, 0.0618280, 0.1791120, 0.1489020, 0.1099720, 0.1978060, 0.1885750, 0.1271390, 0.0360102, 0.0212904, 0.1979290, 0.1803760, 0.1949050, 0.2822160, 0.3322970, 0.1286330, 0.1134640, 0.0358589, 0.0035609, 0.0002349, -0.0072390, -0.0078128, -0.0155750, 0.1212280, -0.0155565, -0.1733020, -0.2342740, -0.1281140, -0.1467340, -0.0712866, 0.0794074, 0.1303980, -0.1982960, 0.0360576, -0.0448275, 0.1662080, 0.1384020, 0.1326770, 0.1459170, 0.3029350, 0.3252320, 0.2184060, 0.2385250, 0.2093870, 0.0815078, 0.0193821, 0.0005960, -0.0001032, 0.0004622, 0.0048623, 0.0029386, 0.1990520, 0.0512813, -0.1613380, -0.2459500, -0.0487823, -0.0668548, -0.1321950, -0.2398020, 0.0190917, 0.1597320, 0.0180978, -0.1801700, 0.0146256, -0.0386617, 0.1078240, 0.1388400, 0.3039140, 0.2627880, 0.1295340, 0.2456630, 0.1991560, 0.0397481, -0.0041773, 0.0000443, 0.0003340, -0.0001067, 0.0003267, -0.0068776, 0.0869925, 0.0559332, -0.0661052, -0.1793070, -0.0390942, 0.0799521, -0.0785479, -0.2969440, -0.2162430, -0.1926300, -0.2686800, -0.2757140, -0.1448420, -0.1568850, 0.0495832, 0.0510182, 0.2425750, 0.1650340, 0.0166180, 0.1739760, 0.1117230, 0.0374263, -0.0053658, -0.0001559, 0.0002804, 0.0001589, -0.0014904, -0.0053577, -0.0775872, -0.0763639, -0.1001690, -0.2108940, -0.2418770, -0.1360660, -0.0842182, -0.2809840, -0.2834330, -0.3393160, -0.3538380, -0.2657010, -0.2551370, -0.1802330, -0.1470820, -0.0071256, 0.1457050, 0.0335622, 0.1368830, 0.1290970, 0.0899891, 0.0131745, 0.0009508, 0.0005985, 0.0001725, -0.0003589, -0.0004953, -0.0205250, -0.0246356, -0.1131690, -0.0526269, -0.1066210, -0.1254200, -0.0935822, -0.0327922, -0.2121350, -0.2446090, -0.3250000, -0.2836540, -0.2056990, -0.1774080, -0.1448780, -0.0530571, 0.0475191, 0.0723412, 0.0720838, 0.0807569, 0.0740009, 0.0450584, 0.0165222, 0.0008558, 0.0005558, 0.0001647, 0.0001110, -0.0002016, -0.0094184, -0.0305125, -0.0180791, 0.0263059, -0.0031151, -0.0167225, -0.1366700, -0.1215650, -0.0280213, -0.0209368, 0.0340788, -0.0063503, -0.0717741, 0.0504475, -0.0423237, -0.0876024, -0.0430445, 0.0529905, 0.0221699, -0.0044425, 0.0122162, 0.0024704, 0.0009162, 0.0010302, -0.0003144, -0.0002559, 0.0000912, -0.0000076, -0.0002897, 0.0177118, 0.0754122, 0.1148810, 0.0893549, 0.0573574, 0.0008010, 0.0098391, 0.0384946, 0.0469515, -0.0561420, 0.0494206, 0.0484990, 0.0422194, -0.0384588, 0.0039983, 0.0052778, 0.0506672, 0.0477501, 0.0119807, 0.0041735, 0.0021210, -0.0001432, 0.0003826, 0.0004688, -0.0003077, 0.0003837, 0.0004590, -0.0001031, 0.0002492, 0.0002781, 0.0019246, 0.0121696, 0.0114597, 0.0030397, 0.0045532, 0.0128841, 0.0173310, 0.0003143, 0.0353379, 0.0385413, 0.0141272, 0.0106257, 0.0399432, 0.0014726, -0.0011148, -0.0036883, 0.0054612, -0.0020025, -0.0000875, -0.0000242, -0.0000991, -0.0004918, -0.0008829, 0.0002879, -0.0001239, 0.0000402, -0.0001279, -0.0002425, -0.0001764, -0.0001847, -0.0005257, 0.0000703, -0.0007776, -0.0004168, -0.0002128, 0.0000677, 0.0001862, -0.0000428, 0.0002512, -0.0006563, -0.0001393, 0.0000207, 0.0002044, 0.0001710, 0.0001758, 0.0000685, -0.0000580, 0.0000602, -0.0006605, -0.0006458, 0.0005823, 0.0002955, -0.0003358, -0.0006827, 0.0000799, -0.0006609, 0.0008380, 0.0024321, 0.0036979, 0.0034917, 0.0069707, 0.0064625, 0.0069134, 0.0113364, 0.0047902, 0.0006575, 0.0029441, 0.0021841, 0.0009232, 0.0011665, 0.0000354, -0.0000429, 0.0008303, 0.0002232, -0.0001196, -0.0001594, -0.0003509, 0.0002589, -0.0006245, 0.0001511, 0.0000990, 0.0007351, 0.0004278, 0.0003731, -0.0000288, 0.0092145, 0.0213731, 0.0246798, 0.0346236, 0.0551576, 0.0812618, 0.0741255, 0.0841423, -0.0036480, -0.0025717, 0.0662287, 0.0756115, 0.0143741, 0.0207043, 0.0177011, 0.0104271, 0.0031636, 0.0009406, -0.0002747, -0.0001070, 0.0000003, -0.0001960, -0.0007699, -0.0030412, -0.0000438, 0.0002916, 0.0047454, 0.0187044, 0.0142107, 0.0716989, 0.0863350, 0.1127550, 0.1628330, 0.1334260, 0.1586940, 0.1281220, 0.1116770, 0.1695030, 0.1469410, 0.1828520, 0.0307743, -0.0451511, 0.0262630, -0.0003869, 0.0161479, 0.0183104, -0.0009636, 0.0055234, 0.0000722, 0.0005106, -0.0002831, -0.0106386, -0.0030221, 0.0042252, 0.0027343, 0.0053442, 0.0693632, 0.1506310, 0.2024280, 0.2071290, 0.1988230, 0.1373730, 0.0434488, 0.0365664, 0.0847576, 0.3220710, 0.2355240, 0.1439780, -0.0253865, -0.1183410, 0.0026178, -0.0082711, -0.0340126, 0.0229903, 0.0325406, 0.0349985, 0.0153425, -0.0002184, -0.0002056, -0.0004693, -0.0029704, -0.0104691, -0.0509274, -0.0215040, 0.0156244, -0.1834860, -0.1243350, 0.0210826, 0.1673100, 0.0915549, -0.0867059, 0.0944918, -0.0301299, 0.2667380, 0.3692990, 0.2898380, 0.3563730, 0.2301430, 0.1350770, 0.0091198, -0.0703843, 0.0421031, 0.1381090, 0.0766670, 0.0167292, 0.0000244, 0.0000944, 0.0014081, -0.0110447, -0.0604362, -0.1293520, -0.1257540, -0.0764200, -0.0807557, 0.0417257, 0.0756927, -0.0028506, 0.0348913, -0.1251180, -0.1026440, 0.0678815, 0.0617004, 0.0200016, -0.0034682, 0.1836880, 0.1647230, -0.0695461, -0.0228227, 0.1226280, 0.0891656, 0.1310060, 0.0296149, 0.0251093, 0.0000162, 0.0050458, -0.0104351, -0.0400122, -0.0476310, -0.0069019, -0.1949530, -0.0131218, 0.0933738, -0.0397615, 0.1111690, 0.1007760, -0.0896285, -0.0735234, 0.1270900, 0.0829104, 0.0020719, -0.2136590, 0.0839038, -0.0977361, 0.0069622, -0.0026042, 0.1703840, 0.1624580, -0.0544764, -0.0901068, -0.0530422, 0.0165433, 0.0000211, -0.0039947, -0.0270556, -0.0114829, 0.0432404, -0.0535555, -0.1010070, -0.0093507, -0.1144030, -0.0967817, -0.0405598, 0.1473320, 0.0284020, 0.1588330, -0.0092920, -0.1188400, 0.1229000, 0.0205746, 0.0607767, 0.2408820, -0.0328506, 0.1533120, 0.1163640, 0.0611872, -0.1069720, -0.0472276, 0.0652693, 0.0087103, -0.0001034, -0.0053511, -0.0152750, -0.0319090, 0.0328559, -0.0037143, -0.0134713, 0.0532460, 0.0297571, 0.0243145, -0.0982942, 0.0130015, -0.1495280, -0.1508030, -0.0579057, -0.0686733, 0.1311720, 0.0449872, -0.0986331, 0.0486785, 0.0582424, 0.0110151, -0.0031025, 0.1858330, 0.1262060, 0.1427040, 0.0460931, -0.0927631, -0.0002072, -0.0058116, -0.0281760, -0.0299237, 0.0361321, -0.0644208, -0.0059588, 0.0668189, 0.1504970, -0.0137682, 0.0989725, 0.0752612, -0.1796440, -0.2513730, -0.0912897, -0.2420770, -0.1988270, -0.0263585, 0.2160240, -0.0904783, 0.1489150, 0.1079770, 0.1196590, 0.2743570, 0.2145360, -0.0454362, -0.0124196, -0.0226879, -0.0002801, -0.0057883, -0.0381934, 0.0044254, 0.1319970, 0.0894876, 0.0498797, -0.0795672, -0.0656142, 0.1231590, 0.0168373, -0.0913151, -0.1126110, -0.0617835, -0.3377050, -0.6030910, -0.5282850, -0.3376000, -0.1494460, -0.0379302, -0.0657298, 0.0315592, -0.0136521, 0.2774610, 0.2286810, 0.0762445, 0.0591841, -0.0015869, -0.0001483, -0.0032717, -0.0147428, 0.0411448, 0.0910228, 0.1592690, -0.0076468, -0.1816590, -0.0544635, -0.0211913, -0.1789510, -0.0068921, 0.0502196, 0.0089416, -0.0736562, -0.4059110, -0.3941470, -0.1997050, -0.4172440, -0.0461468, -0.1663150, 0.0884382, 0.1132190, 0.2321880, 0.1723830, 0.0765465, 0.0216690, -0.0097224, 0.0006374, 0.0001447, -0.0037464, 0.0488364, 0.0153198, 0.2166970, 0.0629692, -0.0929115, 0.0111236, 0.0194151, -0.2701260, 0.1138610, 0.0752817, -0.0102667, -0.0090020, -0.0278465, -0.2746910, -0.3153350, -0.1692310, -0.0128927, -0.0142893, 0.0840565, 0.2323160, 0.1031200, 0.0349007, 0.0574682, 0.0383909, 0.0032595, -0.0001358, 0.0000239, -0.0018432, 0.0002848, -0.1214830, 0.0076322, 0.0699898, -0.1386380, -0.1103190, -0.1480810, -0.1648930, 0.2205050, -0.0546427, -0.0646834, 0.0521876, 0.0116884, -0.3419550, -0.3309180, -0.1982920, -0.2529170, -0.2669460, 0.0529369, -0.1377160, -0.1170240, 0.0455288, 0.0469318, 0.0154435, -0.0001601, 0.0000704, -0.0003215, -0.0027928, -0.0723036, -0.2283590, -0.1422620, -0.1501830, 0.0290210, 0.0518075, 0.0691279, -0.1045890, 0.1311820, 0.0238980, -0.0769533, 0.1989440, -0.1962400, -0.1823050, -0.2650220, -0.0808540, -0.1025650, -0.0768572, -0.1063780, -0.0462250, 0.0980012, 0.1743870, 0.0390697, -0.0068370, -0.0003075, -0.0008530, -0.0002036, 0.0020651, -0.0586077, -0.2959130, -0.2104980, -0.3804220, -0.1766570, -0.1641350, 0.0328936, 0.0865788, 0.1487240, -0.0008368, 0.0669379, 0.0198641, -0.2273910, -0.1981040, -0.3879670, -0.2212160, -0.0346642, -0.1602480, -0.1533590, 0.1109970, 0.2385240, 0.1710940, 0.0601248, 0.0382230, 0.0001785, 0.0000480, -0.0008072, 0.0005905, -0.0221014, -0.2096190, -0.2783250, -0.3371220, -0.1724770, -0.1357850, 0.0363669, 0.2109150, 0.0856303, 0.0346077, 0.1192090, -0.0193874, -0.3681810, -0.3751160, -0.1892340, -0.1787090, 0.0835079, 0.0396159, -0.0163317, 0.0741655, 0.0868667, -0.0215186, -0.0759232, -0.0326678, 0.0028060, -0.0002931, -0.0000261, 0.0050357, 0.0121856, -0.2090750, -0.2117740, -0.1901090, -0.2249820, -0.2146780, -0.0570600, -0.1439650, -0.0588527, 0.0234109, -0.2868820, -0.5589030, -0.4651110, -0.3015450, -0.1517580, -0.0100132, 0.0763687, 0.0179382, 0.0237825, 0.0976861, 0.0758487, -0.0130193, -0.0372305, -0.0321022, -0.0039859, 0.0000219, -0.0001710, 0.0083505, 0.0338994, -0.0999857, -0.0322727, 0.0308061, -0.0220348, -0.0917362, -0.2419690, -0.3486950, -0.3603370, -0.2759240, -0.3217010, -0.5156550, -0.2128380, 0.0387939, 0.2908760, 0.3069530, 0.0946352, 0.0374454, 0.0161458, 0.1000120, 0.1472170, -0.0147218, -0.0143052, -0.0052132, -0.0023328, -0.0002258, 0.0009885, 0.0055305, 0.0590534, 0.0743483, 0.2038000, 0.2374920, 0.1341210, -0.0150296, 0.0281173, -0.1839080, -0.0958355, 0.0763532, 0.2148470, 0.2721940, 0.5529270, 0.3985500, 0.4536390, 0.3219170, 0.2288710, 0.4204930, 0.2869490, 0.2200320, 0.2099390, -0.0080512, -0.0152549, -0.0058347, 0.0002097, 0.0000344, -0.0002595, 0.0012984, 0.0755653, 0.1731970, 0.2322380, 0.3233800, 0.3146340, 0.3775690, 0.3039770, 0.2734070, 0.4893550, 0.2856260, 0.6641730, 0.7800120, 0.6513090, 0.5048650, 0.8235370, 0.4612960, 0.3874430, 0.4250320, 0.1817500, 0.2543120, 0.1953820, 0.0200042, -0.0068580, 0.0000238, 0.0002093, 0.0005247, -0.0000567, 0.0087345, 0.0710000, 0.0814338, 0.1827460, 0.2146200, 0.3578990, 0.4267150, 0.6173130, 0.4396540, 0.6425560, 0.4805030, 0.5287260, 0.2641610, 0.2845300, 0.3553710, 0.4763660, 0.3126790, 0.2132760, 0.1180260, 0.1755110, 0.1453140, 0.1666070, -0.0119575, 0.0010246, -0.0015746, -0.0004656, 0.0000881, -0.0001462, 0.0099507, 0.0543253, 0.0333364, -0.0151951, -0.1219870, 0.0410470, 0.0983564, 0.1502370, 0.1702020, 0.2130100, 0.0586835, 0.2756130, 0.0745355, 0.2117000, 0.1880250, 0.1151040, 0.3428960, 0.2329150, 0.1484300, 0.0800978, 0.1259680, 0.1059750, -0.0169726, 0.0006841, -0.0027393, -0.0001273, -0.0000197, 0.0002155, -0.0054365, 0.0175536, -0.0137220, -0.1145610, 0.0251889, 0.0591579, 0.1147540, 0.0894887, 0.1853030, 0.1908250, 0.3129110, 0.3068510, 0.2497120, 0.2525750, 0.3161450, 0.0486753, 0.2383240, 0.1275910, -0.0436044, -0.0479771, 0.0572824, 0.0219489, 0.0228923, 0.0108112, -0.0002532, -0.0002512, -0.0001445, 0.0002352, -0.0000465, -0.0140354, -0.0694462, -0.0570249, 0.1284200, 0.1502470, 0.1591160, 0.1390940, 0.2369670, 0.0337283, 0.1805700, 0.2456930, 0.1934170, 0.2727720, 0.3138730, 0.1779340, 0.0619430, 0.1566110, -0.0299926, -0.0414530, 0.0129476, -0.0090300, 0.0018660, -0.0015424, 0.0003043, 0.0002041, 0.0001894, 0.0002157, 0.0002543, -0.0001792, -0.0018395, -0.0113745, -0.0268374, -0.0408011, -0.0235955, -0.1369580, -0.0882784, 0.0129199, 0.0761123, 0.0762139, -0.0122165, 0.0014605, 0.0827881, 0.0887761, 0.0025253, -0.0501731, -0.0695284, -0.0499857, -0.0015018, 0.0008505, -0.0001212, -0.0000068, -0.0001827, -0.0000542, -0.0002444, 0.0002974, -0.0004150, -0.0001561, 0.0002273, -0.0005062, -0.0007965, -0.0013520, -0.0027209, -0.0041540, -0.0118698, -0.0039006, -0.0027714, -0.0086517, -0.0103757, -0.0102130, -0.0138188, -0.0169497, -0.0437155, -0.0202168, -0.0319164, -0.0197442, -0.0107832, -0.0032316, -0.0001447, -0.0004819, 0.0000584, 0.0003424, 0.0000382, 0.0000354, -0.0000381, 0.0001100, -0.0002394, -0.0002109, 0.0005580, -0.0003397, -0.0002058, 0.0003787, 0.0001030, 0.0001050, 0.0007080, 0.0001905, -0.0006492, 0.0005332, -0.0002751, -0.0000960, 0.0001052, -0.0001943, -0.0005070, -0.0001592, 0.0005312, 0.0000465, -0.0008165, 0.0004509, 0.0000961, -0.0000156, 0.0009739, 0.0000255, -0.0001374, 0.0001150, -0.0003440, -0.0002131, 0.0001146, 0.0007263, 0.0002338, -0.0001849, -0.0009321, 0.0002371, -0.0000102, 0.0003727, -0.0107735, -0.0284662, 0.0006352, 0.0008861, -0.0018789, -0.0017728, -0.0018896, -0.0000360, -0.0004031, 0.0001006, -0.0003215, 0.0002230, -0.0003548, 0.0001828, 0.0003453, 0.0000681, -0.0004041, -0.0003883, 0.0002593, -0.0002282, 0.0000856, -0.0009316, 0.0029725, 0.0099955, 0.0053114, 0.0098308, 0.0149941, -0.0221268, -0.0198533, -0.0693720, -0.0248028, 0.0053900, -0.0246474, -0.0220958, -0.0169880, -0.0115401, -0.0063783, -0.0027357, -0.0003834, 0.0003028, 0.0004890, 0.0004746, -0.0000520, 0.0005102, -0.0002038, -0.0003640, -0.0023889, 0.0029675, 0.0042933, 0.0046004, 0.0038334, -0.0014835, 0.0031551, 0.0601526, -0.0206106, -0.0674568, 0.0646742, 0.1038370, 0.0637179, -0.0453707, -0.1351290, -0.0684846, 0.0046893, 0.0333727, -0.0189646, -0.0185065, -0.0072713, -0.0005883, -0.0005998, -0.0002058, 0.0001071, 0.0005386, -0.0025711, -0.0015276, -0.0047811, -0.0049099, 0.0032825, -0.0201388, -0.0516258, 0.0110588, 0.0064398, -0.0946092, -0.0618822, 0.0554182, 0.0630299, 0.0187752, 0.0664719, 0.0067097, -0.0991208, -0.0011732, -0.0602682, 0.0117311, -0.0264735, -0.0332011, 0.0371530, 0.0196873, -0.0062889, 0.0013186, 0.0001559, -0.0000137, -0.0008710, -0.0029370, 0.0037094, -0.0017872, -0.0194207, -0.0215687, -0.0370973, -0.0814887, -0.0667282, -0.0536449, 0.0016252, -0.2767920, -0.0970490, -0.1231020, -0.0568555, -0.1031660, -0.2388420, -0.1561500, -0.0840638, -0.0320880, -0.0356110, 0.0093806, -0.0183170, -0.0269313, -0.0049483, 0.0031971, -0.0001500, -0.0001310, -0.0000283, 0.0052497, 0.0445501, 0.1132840, 0.0292447, -0.0714656, -0.1284990, -0.1405130, -0.3562210, -0.2607060, -0.3629900, -0.2143630, -0.2642050, -0.4489730, -0.2875440, -0.3998880, -0.4287510, -0.1873120, -0.1945880, -0.1299300, 0.0514974, 0.1065570, 0.0764092, -0.0185257, -0.0017509, 0.0009962, -0.0000369, 0.0009395, 0.0020438, 0.0160193, 0.0456056, 0.1752780, 0.0880662, 0.0730153, -0.0211587, -0.1558050, -0.2733930, -0.3063070, -0.4169540, -0.2419740, -0.5270970, -0.6494280, -0.7920620, -0.4123130, -0.5274090, -0.2422640, -0.2507320, -0.1382340, -0.1072470, 0.0392851, 0.1526330, 0.0510364, 0.0196848, 0.0001723, 0.0038395, -0.0003645, -0.0026287, 0.0032893, 0.0722722, 0.1838250, 0.1132930, 0.0547493, -0.1861890, -0.1107370, -0.2492620, -0.2681300, -0.4636100, -0.5479150, -0.6150350, -0.5001400, -0.5905500, -0.2881380, -0.1381280, -0.0887129, 0.0824020, 0.0877017, -0.0543956, 0.0196685, 0.1122640, 0.0429678, -0.0057247, -0.0025946, 0.0000947, -0.0006576, 0.0006445, -0.0269732, 0.0173205, 0.1763830, -0.0674269, -0.0737212, -0.1629560, -0.2799820, -0.4531060, 0.0422001, -0.0222150, -0.1550270, -0.3264780, -0.2647420, 0.1326510, 0.1028890, 0.0972796, -0.1164210, 0.0924815, 0.0861632, 0.0020583, 0.1119450, 0.0534937, 0.0013723, -0.0006964, 0.0153000, -0.0005317, -0.0016528, 0.0019511, -0.0372982, 0.0305311, 0.0751802, -0.2645370, -0.0439807, -0.1386770, -0.0594390, -0.0063603, 0.2404580, 0.2436840, 0.0413375, 0.2224430, 0.5841450, 0.2461740, 0.2833400, 0.0225692, -0.1596880, -0.1398960, -0.0473944, 0.1324060, -0.0864396, -0.0171666, 0.0204283, 0.0123603, 0.0042265, 0.0004032, 0.0013631, -0.0054462, 0.0146741, -0.0668903, 0.0931032, -0.1287410, -0.0784006, 0.1588890, 0.2920440, 0.1999240, 0.0687070, 0.2908400, 0.0768390, 0.3360920, 0.3637250, 0.2344410, 0.0379869, -0.0416985, 0.0229010, 0.0250508, -0.0092145, -0.0148793, -0.0474989, -0.0670900, 0.0239305, 0.0036201, -0.0000111, 0.0003750, -0.0005461, -0.0051592, 0.0251107, -0.1746160, 0.0805285, -0.0121027, 0.0355991, 0.3190900, 0.1172050, 0.2689460, 0.1526710, 0.4644770, 0.2405270, -0.0399016, -0.0071819, -0.0396668, 0.0161922, 0.0191002, 0.1180770, 0.2606610, -0.0093761, -0.0064167, -0.0264176, 0.0761461, 0.0484546, -0.0150032, -0.0003721, -0.0002165, 0.0001784, -0.0009571, 0.0538468, -0.0244067, 0.1429060, 0.1474200, 0.0613281, 0.1134820, 0.2452110, 0.1203170, 0.4068060, 0.4396510, 0.0368600, -0.2605920, -0.0195699, 0.1909330, 0.1996170, 0.3028570, 0.1488460, 0.1794400, 0.2024000, 0.2113200, 0.1490450, 0.1186640, 0.0728243, 0.0154776, 0.0004825, 0.0000408, -0.0008000, -0.0000983, 0.0707284, 0.0943884, 0.1912730, 0.0192308, 0.1176890, 0.1749150, 0.3184200, 0.2048690, 0.3336100, 0.2800250, -0.2198310, -0.1068730, 0.0650950, 0.2450160, 0.2453370, 0.0977683, 0.2262150, -0.0282979, 0.1412980, 0.1827180, 0.1401480, 0.1096750, 0.0310137, 0.0142435, -0.0002802, -0.0002303, 0.0004748, 0.0068242, 0.0751391, 0.1297940, 0.2207560, 0.0699316, -0.0523980, -0.0443265, 0.2769900, 0.1019100, 0.1508960, 0.0041877, -0.1655250, -0.0531728, 0.1779840, 0.1989950, 0.1459290, 0.0704541, 0.2839490, 0.1262960, 0.1591920, 0.1147040, 0.1176160, 0.0760686, 0.0518918, 0.0720101, 0.0016305, -0.0000515, -0.0001445, 0.0111019, 0.0596546, 0.0239335, 0.1808610, 0.1828290, 0.1981340, 0.2329360, 0.1422650, -0.0588794, -0.0212451, -0.0063478, 0.0513011, 0.1512050, 0.4961230, 0.2524570, 0.2612900, 0.3378830, 0.3043320, 0.2605880, 0.3355750, 0.0735907, 0.1898040, 0.0854379, 0.0719744, 0.0543447, 0.0034687, -0.0004741, 0.0002844, 0.0369999, 0.0442790, 0.0624468, 0.1661920, 0.2196100, 0.1965290, 0.2433180, 0.1776280, -0.1840530, -0.1200820, -0.0986597, 0.1689960, 0.1227920, 0.0814610, 0.2266090, 0.1635210, 0.3397650, 0.0798064, 0.1859550, 0.4355450, 0.2380950, 0.1657020, 0.0459649, 0.0064484, 0.0089797, 0.0053531, -0.0011367, -0.0002771, 0.0187713, 0.0687771, 0.1708560, 0.1556230, 0.1227030, 0.0340230, 0.0078842, -0.0943750, -0.3851510, -0.1395030, 0.1696830, 0.2350200, 0.1630380, 0.0555301, 0.2122040, 0.1473530, 0.1516320, -0.0383342, -0.0053052, 0.1742360, 0.1567270, 0.1621280, 0.0263881, -0.0226242, -0.0036312, 0.0018674, -0.0005091, -0.0013120, 0.0073003, 0.0876729, 0.1604510, 0.2476600, 0.0470095, -0.0393842, -0.0857710, -0.0520669, -0.0740763, -0.0154387, -0.0800177, 0.2823130, 0.3633270, 0.2512750, 0.2391360, 0.0716861, -0.0444007, -0.3665010, -0.0974556, -0.0465821, 0.0311561, 0.0353773, -0.0604992, -0.0300282, 0.0129890, -0.0003363, 0.0000497, -0.0009274, 0.0172280, 0.0554337, 0.0336347, 0.0502999, -0.0436681, 0.1121800, 0.0311693, -0.0786873, -0.0290120, 0.1204600, 0.0997871, 0.2148610, 0.0269280, -0.0020461, 0.0427271, -0.1555860, -0.1647280, -0.4857320, -0.1512940, -0.1988570, -0.0862612, -0.0132181, -0.1338830, -0.0505692, 0.0035393, 0.0002477, 0.0001846, 0.0002565, 0.0276484, 0.0597519, 0.0280230, -0.0147549, -0.1714800, -0.0830978, 0.0457314, 0.0042722, -0.0846768, 0.0700133, -0.0338396, -0.1990260, -0.3800180, -0.1680570, -0.1033700, -0.0083295, -0.2495280, -0.2674240, -0.3033490, -0.2809050, -0.1005140, -0.1097650, -0.1361360, -0.0098641, 0.0023213, 0.0001104, 0.0000045, 0.0002821, 0.0033057, -0.0109433, 0.0051239, -0.0859602, -0.1980400, -0.1572150, -0.1774130, -0.1223470, -0.1177300, -0.1461550, -0.2484330, -0.2252530, -0.3728080, -0.1380510, -0.0480899, -0.1537300, -0.1502650, 0.0861211, -0.1440680, 0.0276722, -0.0831270, -0.1735370, -0.1349790, 0.0103089, 0.0091173, 0.0000212, -0.0003265, 0.0002147, 0.0003273, -0.0074792, -0.0024645, -0.1042890, -0.1807950, -0.1881680, -0.2120980, -0.1387240, -0.0573749, -0.1509450, -0.1119540, -0.2427960, -0.0330267, -0.2780910, -0.3884500, -0.1941210, -0.0942919, -0.0359680, -0.1487830, 0.0119438, -0.1773490, -0.2022660, -0.1597380, 0.0139725, 0.0094393, -0.0005161, 0.0000369, -0.0005402, -0.0000464, 0.0048620, -0.0079141, -0.0775069, -0.0815632, -0.2062380, -0.2323140, -0.2066790, -0.2247990, -0.1367860, -0.3112730, -0.1158950, -0.0663380, -0.3148830, -0.0586322, -0.0686283, -0.0913629, -0.0434077, -0.1349810, 0.0855351, -0.0596009, -0.1134020, -0.0414042, 0.0021231, -0.0006090, 0.0000423, -0.0001679, 0.0000074, -0.0001975, 0.0014532, -0.0058167, -0.0598531, -0.0497403, -0.1316710, -0.3173730, -0.3076360, -0.1809830, -0.2251200, -0.2747790, -0.2171200, -0.3051800, -0.2404630, -0.2684190, -0.1822010, -0.1346460, -0.3647050, -0.2186310, -0.1234990, -0.0327516, -0.0019696, -0.0008527, -0.0006432, 0.0004424, 0.0003079, 0.0005003, 0.0002792, -0.0000427, 0.0000708, -0.0071151, -0.0420384, -0.0569232, -0.0604198, -0.0986802, -0.1424240, -0.1922580, -0.2522990, -0.1906630, -0.2554670, -0.4489940, -0.3303660, -0.2790140, -0.2451750, -0.1938310, -0.1526330, -0.1703070, -0.1322330, -0.0287627, -0.0086620, -0.0004605, -0.0000598, -0.0003173, 0.0004521, -0.0001761, -0.0002852, 0.0003095, 0.0001875, 0.0004268, 0.0011309, 0.0000556, -0.0002780, 0.0003812, 0.0018756, 0.0006273, -0.0043383, 0.0004548, -0.0006687, -0.0535198, -0.0368489, -0.0216304, -0.0105858, -0.0360878, -0.0112738, -0.0193764, -0.0160202, -0.0056689, 0.0002552, 0.0007161, -0.0001814, 0.0000232, 0.0002708, 0.0003551, 0.0005187, 0.0003020, 0.0003328, -0.0001752, -0.0004018, 0.0003139, -0.0001141, -0.0000594, -0.0006480, -0.0002238, -0.0000147, -0.0005517, 0.0002423, -0.0003348, -0.0001364, 0.0002494, 0.0001533, 0.0002993, 0.0004265, 0.0003187, 0.0004052, 0.0001739, 0.0002136, -0.0002948, 0.0000116, 0.0002932, 0.0001363, -0.0000620, 0.0003657, 0.0003729, -0.0003096, 0.0002717, -0.0004565, 0.0112228, 0.0183403, 0.0235827, 0.0057687, 0.0031560, 0.0032380, 0.0072420, 0.0143323, 0.0093686, 0.0041376, 0.0110916, 0.0053898, 0.0001885, 0.0010603, -0.0000639, 0.0003452, 0.0032317, 0.0053160, 0.0002847, 0.0000500, 0.0001512, 0.0003906, -0.0000076, 0.0001705, 0.0005413, 0.0001568, 0.0001892, 0.0004514, 0.0080996, 0.0343531, 0.0391602, 0.0235996, 0.0302061, 0.0314089, 0.0474197, 0.0675709, 0.0613952, 0.0105826, 0.0091882, -0.0260070, -0.0202133, -0.0157087, -0.0062538, 0.0001233, 0.0029874, 0.0034398, -0.0000410, 0.0001368, -0.0005295, 0.0002186, -0.0002573, 0.0006984, -0.0001339, 0.0003205, -0.0005957, -0.0003716, 0.0507030, 0.0708823, 0.0457716, 0.0660915, 0.0586532, 0.0377397, 0.0320708, 0.1511950, 0.1080030, 0.0484198, -0.0047176, -0.0543424, -0.0304982, 0.0009859, -0.0030088, -0.0189751, -0.0199991, 0.0068705, 0.0049668, -0.0000801, 0.0008012, 0.0001350, -0.0000430, -0.0002396, -0.0002718, -0.0015823, -0.0027852, -0.0062460, 0.0576299, 0.0712897, 0.1073420, 0.1933330, 0.1173550, 0.0754353, 0.1771950, 0.2865300, 0.3207680, 0.2184270, 0.1331650, 0.1392510, -0.0332170, -0.1015830, 0.0076797, -0.1110290, -0.0519520, -0.0412496, -0.0122369, 0.0465389, 0.0325486, 0.0056600, -0.0000985, 0.0002646, 0.0000096, 0.0012641, 0.0322431, -0.0199929, 0.0536915, -0.0243683, -0.1506250, -0.1843920, 0.0775362, 0.0983231, 0.0187073, 0.2026660, 0.1036410, 0.0922238, 0.0672866, 0.1376690, 0.1634560, 0.1593850, 0.2029650, 0.1346780, 0.0889407, -0.0312115, -0.0189451, 0.0704145, 0.0417164, 0.0035033, 0.0003592, 0.0002949, -0.0109323, -0.0213377, -0.0170167, -0.0866186, 0.0007698, -0.0345805, -0.1727860, -0.1015200, 0.0679172, -0.1926950, 0.0580117, -0.0584742, -0.0932499, 0.0823743, -0.1259490, -0.1553810, -0.0030093, 0.0335574, -0.0772939, -0.0587690, 0.0573593, 0.0689531, 0.0214623, 0.0941677, -0.0206952, -0.0001135, 0.0002220, -0.0003453, -0.0143362, -0.0825675, -0.0141878, 0.1753560, 0.0937152, 0.0175125, 0.0646582, -0.1485390, -0.1326710, 0.0040134, 0.0696659, -0.0873961, 0.0296949, 0.3152010, 0.0821108, -0.0727521, 0.1921850, 0.0930965, 0.0369348, -0.0634680, 0.0635810, -0.0085369, -0.0790158, 0.0400938, -0.0850599, -0.0009624, 0.0001397, -0.0043500, -0.0196431, -0.0694905, -0.0392903, -0.0174423, 0.0584353, 0.0243914, -0.0699589, 0.0186415, 0.1406960, -0.0343031, -0.0265320, 0.1011440, 0.0495865, -0.0357401, 0.1197510, -0.0822424, -0.0659674, 0.0424991, 0.1341010, -0.0248103, -0.0229683, 0.0993981, -0.0760581, 0.0234603, 0.0603935, 0.0077420, 0.0000161, -0.0077670, -0.0210139, -0.0784834, -0.1517470, 0.0132167, -0.0468820, -0.1020040, -0.1542950, -0.0499794, 0.1228270, -0.0687419, -0.1381870, -0.0469307, -0.2052870, -0.0745665, -0.0381001, -0.3417220, -0.2714490, -0.0114146, -0.1937850, -0.0210956, 0.0629940, 0.2605350, 0.0546518, 0.1362970, 0.0710392, -0.0681784, -0.0002666, -0.0038954, -0.0227492, -0.1439160, -0.1663280, -0.0342440, -0.0481977, 0.0315747, -0.1885280, -0.1697750, 0.0868362, -0.1562750, -0.1232500, -0.0244713, 0.0621352, -0.0604270, -0.1488120, -0.0585787, -0.0549091, -0.1377180, -0.1235980, 0.0208757, 0.1016100, 0.2408370, 0.0879110, -0.1216140, -0.0058592, -0.0127669, -0.0004634, -0.0032116, -0.0301878, -0.0797612, -0.0782468, -0.1175550, -0.0415251, -0.0202611, -0.2440580, -0.1188160, -0.0888533, -0.2606750, 0.0208132, 0.1399230, -0.0888353, -0.0862226, -0.0543292, -0.2732390, -0.0877335, -0.1174510, -0.1509760, -0.1446570, -0.1400610, 0.1389940, 0.1948210, 0.0058136, 0.0398716, 0.0013228, -0.0005355, -0.0027428, -0.0228870, 0.0366554, -0.0199716, 0.1624410, 0.0984326, -0.0307527, -0.1253810, 0.1624980, -0.0945160, 0.0283471, 0.1848140, 0.0631622, -0.1360820, -0.3284210, -0.2890360, -0.2513700, -0.2208420, -0.0743553, -0.1353910, -0.0993422, -0.1281150, 0.1683550, 0.2394970, 0.0228459, -0.0271489, -0.0116436, 0.0001792, -0.0002866, -0.0100131, 0.0694456, -0.1146890, -0.0277410, 0.0386357, -0.1075190, 0.1258710, 0.1524510, -0.0600960, 0.0334671, 0.1836600, 0.0004525, -0.0892102, -0.1484590, -0.0978396, -0.1093180, -0.0571367, -0.0138235, -0.1454350, -0.0558689, 0.0066936, 0.1445100, 0.1472070, 0.0162176, 0.0076069, 0.0054883, 0.0004558, -0.0020305, -0.0059717, 0.0001710, -0.1090370, -0.1633150, 0.0913447, -0.1760230, -0.1646180, -0.1663990, 0.0367390, 0.0214537, -0.0217694, 0.0123639, -0.0466874, -0.1588900, -0.0370062, -0.0773255, -0.1318670, -0.1611710, -0.1416910, -0.1479080, -0.1627090, -0.0548673, 0.1603750, 0.1296680, 0.0502945, 0.0001916, -0.0002165, -0.0050998, 0.0120536, -0.0296345, -0.0647826, -0.1026930, 0.0550306, 0.0490991, 0.0027860, -0.0414431, -0.1837340, -0.1345400, 0.0195469, 0.0910577, -0.0422826, -0.0777945, -0.0858808, -0.3106690, -0.2300440, -0.1604650, -0.2390510, -0.3425970, -0.2503330, -0.0389515, 0.2893690, 0.1902370, 0.0136305, 0.0053194, 0.0003261, -0.0019747, 0.0415917, -0.0004516, 0.0072701, 0.0074013, -0.0196739, -0.0947536, -0.1241380, -0.0954589, -0.0478539, -0.2314890, -0.2596540, -0.1111690, -0.0471048, -0.1516990, -0.0314779, -0.1392140, -0.2133410, -0.0638685, -0.0530178, -0.1364890, 0.0742436, 0.2519280, 0.3038420, 0.1549400, 0.0409658, 0.0034125, -0.0005370, -0.0008240, 0.0442147, 0.0537073, 0.0884668, 0.2020770, 0.2543710, 0.1872840, 0.0920075, -0.0497808, -0.0955173, -0.1995530, -0.1476700, -0.0765771, 0.0420555, -0.1465810, -0.0068802, 0.0481597, -0.1388960, 0.1515910, 0.2032170, 0.0304176, 0.1394120, 0.1098770, 0.1130130, 0.0054299, -0.0201826, 0.0191591, -0.0008107, -0.0001350, 0.0037364, 0.0540816, 0.1479010, 0.4106400, 0.6047710, 0.6365410, 0.6867730, 0.7145780, 0.5474410, 0.2339010, 0.1867860, 0.0623436, 0.1565840, 0.2333230, 0.2385360, 0.1611990, 0.2302480, 0.3566320, 0.2197280, 0.1476000, 0.2734310, 0.2899090, 0.1717250, -0.0022521, -0.0334410, 0.0019383, 0.0002932, -0.0007605, -0.0010681, 0.0055671, 0.1649090, 0.4294460, 0.6287730, 0.7324400, 1.0577900, 1.0020000, 1.0068300, 0.7061640, 0.6463210, 0.4946490, 0.3048910, 0.3286160, 0.3072630, 0.3611470, 0.3069650, 0.2769810, 0.3752320, 0.3572700, 0.4636630, 0.3531960, 0.1434870, -0.0052795, 0.0049304, -0.0005065, 0.0003983, -0.0001744, -0.0059607, -0.0030498, 0.1640460, 0.3308590, 0.3961110, 0.4149530, 0.4681170, 0.4965790, 0.6156330, 0.4343390, 0.5668210, 0.3756740, 0.1040980, 0.1317480, 0.1013580, 0.1428230, 0.0918510, 0.2241340, 0.4127080, 0.2398720, 0.2099930, 0.1619750, 0.0723823, -0.0175096, 0.0019191, -0.0001491, -0.0000457, 0.0002574, -0.0173232, -0.0087444, -0.0088669, 0.1138380, 0.0408292, -0.0133463, -0.0842757, -0.2620400, -0.1342030, 0.0136585, 0.0445652, 0.2167170, 0.1561090, 0.1088770, -0.0554909, 0.2937660, 0.0251319, 0.2101180, 0.2646770, 0.0997591, 0.1547150, 0.0795262, -0.0153148, -0.0064393, 0.0015487, -0.0002741, -0.0002997, -0.0005403, -0.0000312, 0.0142004, -0.0601231, -0.0898230, -0.1865150, -0.2323590, -0.3014690, -0.2677550, -0.3569540, -0.1537100, -0.0022344, 0.1391760, 0.2532640, 0.1284230, 0.1117270, 0.1030270, 0.1998710, 0.2823050, 0.2989400, 0.2969310, 0.1530160, 0.0499829, -0.0400802, -0.0224593, -0.0012018, -0.0002283, -0.0002858, -0.0001591, 0.0038027, -0.0162507, -0.0941307, -0.1661200, -0.3057120, -0.2679230, -0.0002709, 0.1114460, -0.0437642, 0.1276070, 0.2148650, 0.1115490, 0.0413592, 0.3790810, 0.3099640, 0.2263650, 0.2102370, 0.2717230, 0.3138670, 0.2688700, 0.1148860, -0.0082471, -0.0502854, -0.0037002, -0.0009046, -0.0003128, 0.0001568, -0.0005325, 0.0002177, -0.0298670, -0.1207990, -0.2911360, -0.2746200, -0.2096940, -0.0558059, -0.0179778, 0.0373629, 0.0208881, 0.2017060, 0.1064660, 0.2033440, 0.2563860, 0.2183960, 0.1351350, 0.2367830, 0.2440300, 0.1246270, 0.0591720, 0.0180692, -0.0297198, 0.0007912, 0.0087388, 0.0017299, 0.0001969, 0.0001775, -0.0001968, -0.0003132, -0.0122057, -0.0946217, -0.1909330, -0.0413830, -0.0665283, -0.0788102, -0.0668671, 0.0457767, -0.1278320, 0.0111990, -0.0458726, -0.1054960, 0.0135429, -0.0648913, 0.0117382, 0.0391899, 0.0483155, -0.0205338, -0.0219184, -0.0500767, -0.0451488, -0.0112216, 0.0019304, 0.0018123, -0.0000519, -0.0006670, 0.0004739, 0.0001584, 0.0002758, -0.0028934, -0.0217383, -0.0746328, -0.0705920, -0.0331629, -0.0631927, -0.0928006, -0.0113001, -0.0101107, -0.0601898, -0.1776780, -0.1570890, -0.0975332, -0.0222025, -0.0239653, -0.0591875, -0.0417366, -0.0043270, -0.0075527, -0.0010349, -0.0013422, -0.0002497, -0.0007777, -0.0005507, 0.0001248, 0.0001206, 0.0007561, -0.0007554, 0.0000665, -0.0004785, -0.0003000, -0.0004076, -0.0005287, -0.0019365, -0.0067279, -0.0015729, -0.0013919, -0.0051022, -0.0086657, -0.0111046, -0.0112947, -0.0077739, -0.0239337, -0.0221100, -0.0214261, -0.0143807, -0.0124298, -0.0033216, -0.0005487, 0.0003225, -0.0000655, 0.0000878, -0.0002414, 0.0000090, -0.0000226, 0.0000213, 0.0006067, -0.0001511, -0.0002873, -0.0001805, -0.0002754, 0.0001692, -0.0004714, -0.0002087, 0.0002935, 0.0001553, 0.0003969, -0.0001855, -0.0002091, -0.0001612, 0.0003082, 0.0001142, -0.0002632, -0.0001139, 0.0003618, -0.0000635, 0.0001686, 0.0000200, 0.0001194, -0.0012246, -0.0001128, 0.0003264, -0.0002124, 0.0000536, -0.0006731, -0.0002302, 0.0000665, 0.0000588, 0.0001500, 0.0001391, 0.0005027, -0.0001668, -0.0005007, 0.0005176, 0.0001211, 0.0004445, -0.0000392, -0.0005333, -0.0001304, 0.0001232, 0.0000903, -0.0001500, 0.0000722, 0.0001025, -0.0005245, 0.0000485, -0.0001466, 0.0001550, -0.0000406, -0.0001634, 0.0003061, -0.0003499, 0.0002779, -0.0003453, -0.0002117, 0.0005892, -0.0009970, -0.0265259, -0.0068977, -0.0055953, -0.0226376, -0.0064452, 0.0355830, 0.1188330, 0.0543721, 0.0310454, 0.0387853, 0.0259353, 0.0135301, 0.0076428, 0.0076672, 0.0023213, -0.0000386, 0.0005270, 0.0002732, 0.0004826, -0.0005704, 0.0001324, 0.0002956, -0.0013279, -0.0010898, 0.0060073, 0.0043866, -0.0039924, -0.0382105, -0.0939998, -0.1168910, -0.1668870, -0.0243259, -0.0689203, 0.0149166, 0.1514990, 0.1125240, -0.0349999, -0.0033136, -0.0088279, -0.0420158, -0.0581532, -0.0995627, -0.0884342, -0.0329392, -0.0031704, -0.0005167, -0.0001669, -0.0006563, -0.0004955, 0.0014064, 0.0012263, 0.0133217, 0.0240898, 0.0014960, -0.0570309, -0.0442859, -0.1231090, -0.0181724, 0.0938571, 0.0651208, 0.0816190, -0.0992325, 0.2008420, -0.0938417, -0.2266560, 0.0228508, -0.0180299, -0.1690980, 0.0110137, 0.0157944, 0.0297365, 0.0957217, 0.0640032, 0.0114756, -0.0012880, 0.0001114, 0.0001151, 0.0000067, -0.0002879, 0.0302617, 0.0855760, 0.0648066, -0.0153665, -0.1350180, -0.1091850, 0.0029114, 0.0804321, -0.0898388, 0.0933980, -0.0463130, -0.0340629, 0.1160210, -0.0720370, -0.2061830, -0.1034130, 0.0094182, -0.1867990, 0.0385421, 0.1605410, 0.1352520, 0.0606430, -0.0166489, -0.0022776, 0.0000258, -0.0002423, 0.0058787, -0.0358477, -0.0053540, -0.0059985, -0.0366892, -0.0743204, -0.0617858, -0.0674967, -0.0218747, 0.0890424, -0.0441475, 0.1201240, 0.0240974, -0.0333627, 0.0235203, 0.0706685, 0.0490935, 0.0328987, 0.1201450, 0.0725916, 0.0899563, 0.0882353, 0.1690270, 0.0951065, 0.0496011, 0.0057187, 0.0003625, 0.0012500, -0.0146586, -0.0795440, 0.0138955, 0.0247752, -0.0729291, -0.0869075, 0.0398710, -0.1237630, -0.0933422, 0.0830247, -0.0229379, 0.0247987, 0.3158980, -0.0419605, 0.0903054, -0.1309850, 0.0348508, -0.0468858, 0.0372939, 0.0337401, 0.0108507, -0.0004469, 0.1708660, 0.1030710, 0.0275429, 0.0032317, -0.0001292, -0.0034176, -0.0319217, 0.0023515, 0.1047270, 0.0726563, -0.1088210, -0.0800659, 0.0634917, 0.0892951, 0.0331126, 0.0714469, 0.0311240, 0.0856543, -0.0822687, 0.1013160, 0.1286980, 0.0779899, -0.0265762, -0.0955616, -0.0766628, -0.1225740, -0.1514360, -0.0604954, 0.1681720, 0.1613310, 0.0289942, 0.0031998, 0.0002931, -0.0035142, 0.0028366, 0.0330754, 0.1188430, -0.0220464, 0.0281535, 0.1263200, -0.0383448, -0.0285875, 0.0265331, 0.0302431, -0.0253012, 0.0650853, -0.0521222, -0.0225784, -0.2303080, -0.1198450, 0.1491370, -0.0764776, -0.0843875, -0.1068480, 0.0056295, -0.1185100, 0.0717700, 0.1318260, 0.0258278, 0.0002448, -0.0004302, -0.0040803, 0.0043672, 0.0949550, 0.0131015, -0.0480760, 0.0268525, -0.0740909, 0.0358537, -0.2511750, 0.0195998, -0.1195170, -0.0173106, 0.0973157, -0.0997068, -0.1864850, -0.4072540, -0.0623885, -0.0206377, 0.0180846, 0.0770488, 0.0859046, -0.0924351, -0.0739206, 0.0943645, 0.1988070, 0.0617925, 0.0008231, 0.0001205, -0.0045417, -0.0158017, -0.0322928, -0.0134399, -0.0304666, -0.0625784, -0.0975436, -0.1787940, -0.1286710, -0.0044881, -0.1461410, 0.1189790, 0.1600030, -0.0133272, -0.0473433, -0.0414527, -0.0892999, 0.0845173, -0.0171811, 0.0297510, -0.0088761, 0.1094680, 0.0446315, 0.0053838, 0.0654074, 0.0623066, 0.0020281, 0.0007770, -0.0022035, -0.0134720, -0.1077350, -0.0205921, -0.0470017, -0.0133382, 0.0113439, 0.0179050, 0.0494546, 0.0837060, 0.1543680, 0.1862430, 0.2044250, 0.0049696, -0.0757322, -0.1752210, -0.2202580, -0.1409120, -0.3801080, -0.1053250, -0.0289764, -0.0088831, -0.0538387, -0.1428460, -0.0521636, 0.0297966, 0.0012192, -0.0003511, -0.0005391, -0.0172078, -0.1168990, -0.1095610, 0.0574124, -0.0028746, 0.0118378, -0.0635998, -0.0007063, 0.0502710, 0.1213330, 0.0360183, -0.0950098, 0.0945539, -0.1171310, -0.0650232, -0.0825126, -0.1418940, -0.1351640, -0.0622693, -0.1029560, -0.1484510, -0.1083870, -0.0965014, -0.0779612, -0.0030281, -0.0006815, 0.0000055, 0.0045423, -0.0095737, -0.0659344, -0.1024100, -0.1762500, 0.0722422, 0.1443530, 0.1070720, 0.0553983, -0.0850048, -0.1399950, 0.1507950, -0.0122785, 0.1011750, 0.1329700, -0.0964142, -0.1599240, -0.0327079, -0.1823090, -0.0215653, 0.0531714, -0.0435292, 0.0223611, -0.1088960, -0.0840493, -0.0087305, -0.0003295, 0.0002111, 0.0123980, 0.0110879, -0.0625444, -0.1436000, -0.1845400, -0.0880179, -0.1646470, 0.0281089, 0.2006720, 0.4041030, 0.2793220, 0.0355695, -0.0448817, -0.0311491, 0.0265823, -0.0068220, -0.3711510, -0.1272810, -0.0989433, 0.0888140, 0.1460230, 0.0444845, 0.0793581, -0.0461757, -0.0786502, 0.0103338, -0.0004926, -0.0007431, 0.0057323, 0.0248709, -0.0319338, -0.2509840, -0.3166590, -0.5769630, -0.6132210, -0.4615900, -0.1279160, 0.2598070, 0.2849440, 0.4371050, 0.1577410, -0.1093000, -0.0983880, -0.2173100, -0.2517010, 0.1210340, 0.0479598, 0.0174616, -0.1215820, 0.0879858, 0.0189646, 0.0835902, -0.0715620, -0.0285769, -0.0009439, -0.0001857, 0.0025812, 0.0228019, 0.0320375, -0.3223960, -0.5687830, -0.7439900, -0.7265680, -0.8938860, -1.1516100, -0.7410690, -0.4051830, -0.2359980, -0.1867010, -0.1934530, -0.1186680, -0.3184840, 0.0112948, 0.1644790, -0.0119204, 0.0375365, -0.1944510, -0.0781851, 0.0061161, -0.0586507, -0.0507517, -0.0134495, 0.0001577, -0.0006676, -0.0002405, 0.0125999, 0.0721386, -0.1981620, -0.4619450, -0.4260850, -0.5773880, -0.9519720, -1.4328000, -1.4370300, -1.3551800, -1.1509600, -0.8609490, -0.4629940, -0.2456560, 0.1114630, 0.1080810, -0.0144294, 0.0407454, 0.0630749, 0.1095040, 0.0018691, -0.0340927, -0.1294240, -0.0254724, -0.0076610, 0.0004761, -0.0002311, -0.0022570, 0.0094782, 0.1017070, -0.0134275, -0.1548270, -0.1033760, -0.2128880, -0.2396710, -0.3225400, -0.5763520, -0.7475230, -0.5709620, -0.3138520, -0.0403431, 0.1769620, 0.3475730, -0.0967413, 0.1178510, -0.0667710, 0.0781586, 0.0254952, 0.0412074, 0.1770630, -0.0255541, -0.0181189, -0.0042351, 0.0003477, 0.0001544, 0.0012589, -0.0173011, 0.0440337, 0.0375434, 0.0850026, 0.1246240, 0.0745478, 0.2328490, 0.4226520, 0.3194840, 0.2991930, 0.1778940, 0.1382430, 0.1351890, 0.0422190, -0.0608712, 0.1707180, 0.2553230, 0.0580939, 0.1151300, -0.0304242, 0.0574955, 0.0774753, -0.0152857, -0.0150723, -0.0021976, 0.0008154, -0.0003989, 0.0006658, -0.0742579, 0.0352023, 0.1339870, 0.1655110, 0.2986990, 0.2984170, 0.3242840, 0.3210750, 0.3844170, 0.3080600, 0.2961530, 0.2228370, 0.1417550, 0.1732030, 0.0441329, -0.0345810, 0.0452422, 0.0114853, 0.1327890, -0.0674966, -0.0193402, 0.0366451, -0.0386941, -0.0114570, -0.0002988, -0.0005109, -0.0000757, 0.0003058, -0.0621697, 0.0029340, 0.1244440, 0.2369910, 0.1324550, 0.0983666, 0.1431430, -0.0054900, 0.2453560, 0.3387890, 0.2538780, 0.2050660, -0.0437504, 0.1083900, -0.0694665, -0.0538347, -0.0681716, 0.0534489, 0.2764170, -0.0606662, 0.0560743, -0.0021831, -0.0233156, -0.0202624, -0.0018244, 0.0000938, 0.0000849, 0.0005257, 0.0237270, 0.0646798, 0.1800380, 0.3242530, 0.1259350, 0.1238310, 0.2838370, 0.1224960, 0.3287880, 0.2099930, 0.0787873, 0.1790120, 0.1970370, 0.0496227, 0.1620580, 0.1338970, 0.0274498, 0.0620721, 0.0689988, -0.0371711, -0.0341962, -0.0250594, -0.0042410, -0.0176874, -0.0002464, 0.0005810, -0.0001897, -0.0002038, 0.0102114, 0.0496480, 0.1139210, 0.1658440, 0.1913920, 0.3324600, 0.2798500, 0.1129650, 0.2204280, 0.1128100, 0.1425320, 0.1466530, 0.1506340, -0.0466987, -0.1477560, 0.1438040, -0.0455150, -0.1714680, -0.0514845, 0.0332762, 0.0312644, 0.0001127, -0.0101019, -0.0005786, 0.0003212, 0.0000508, 0.0002853, -0.0001765, 0.0011529, -0.0007762, 0.0302447, 0.0945158, 0.0714078, 0.1273480, 0.0904328, 0.1106020, 0.2161820, 0.0907927, 0.1993230, 0.2623830, 0.0416773, 0.0479701, 0.0041274, -0.0083504, 0.0110816, 0.0259763, 0.0338511, 0.0533938, 0.0502915, 0.0038729, 0.0018029, 0.0008949, 0.0002464, -0.0004074, 0.0000083, -0.0004999, 0.0001912, 0.0000172, 0.0032334, 0.0469747, 0.0567533, -0.0010801, -0.0665163, -0.0880507, -0.0249853, 0.0453898, 0.0582845, 0.0296592, -0.0501929, -0.0310104, 0.0551959, 0.0326703, 0.0383817, -0.0105483, 0.0191840, 0.0347063, 0.0053646, 0.0024714, -0.0006870, 0.0006451, 0.0005081, 0.0006234, -0.0007410, 0.0000765, 0.0004497, -0.0003275, -0.0002312, -0.0001814, -0.0005759, -0.0026634, -0.0054587, -0.0111856, -0.0272532, -0.0178789, -0.0177453, -0.0314619, -0.0116301, -0.0077190, -0.0112476, -0.0109298, -0.0098238, -0.0173362, -0.0078273, -0.0052004, -0.0033361, -0.0000578, -0.0005897, -0.0001555, -0.0003009, 0.0001206, -0.0000255, -0.0006214, -0.0001690, 0.0002290, -0.0001226, 0.0004559, 0.0002258, 0.0000357, 0.0006472, -0.0006861, -0.0001086, -0.0000049, 0.0009369, 0.0014487, -0.0006790, 0.0007811, 0.0001963, -0.0001706, -0.0000544, 0.0004220, 0.0002943, 0.0002625, 0.0001314, 0.0000481, -0.0004646, -0.0000098, 0.0006351, -0.0008077, 0.0000064, 0.0004322, -0.0003606, -0.0000366, -0.0001558, -0.0001882, -0.0001293, 0.0006713, 0.0035637, 0.0051734, 0.0084271, -0.0083581, 0.0023687, 0.0127554, 0.0105163, 0.0150053, 0.0044459, 0.0090993, 0.0114365, 0.0059218, 0.0118167, 0.0085972, 0.0040761, 0.0015388, -0.0001192, 0.0002006, 0.0001008, -0.0002503, 0.0001354, 0.0000178, 0.0004244, 0.0003102, 0.0003851, -0.0005625, -0.0014548, 0.0038359, 0.0118860, -0.0034296, 0.0064168, 0.0256739, 0.0461027, 0.0277961, 0.0376227, 0.0727974, 0.0684739, 0.0353942, 0.0414673, 0.0859232, 0.0144759, -0.0028965, 0.0059030, 0.0047823, -0.0009333, -0.0009385, -0.0000076, 0.0004199, -0.0001599, -0.0000552, 0.0000401, 0.0022989, 0.0154457, 0.0569289, 0.0609768, 0.0666180, 0.0843029, -0.0004106, -0.0151033, -0.0321743, 0.1021310, 0.1429760, 0.1324550, 0.1426090, 0.0090150, -0.0497590, 0.0378625, 0.1001390, 0.0663022, -0.0134753, -0.0289045, -0.0055842, 0.0139446, 0.0002855, 0.0003689, 0.0001227, 0.0000122, -0.0003094, -0.0001131, 0.0048212, 0.0142558, 0.0464433, -0.0063299, 0.0178399, 0.0840402, 0.0136487, 0.1181830, -0.0223144, 0.0585246, -0.0890620, -0.1976770, 0.0116159, -0.0390407, 0.0041239, 0.1107390, 0.0630186, 0.0796663, 0.2144410, 0.1166020, 0.0101508, -0.0057929, -0.0029185, 0.0002436, 0.0005036, 0.0003833, 0.0001179, -0.0011629, 0.0165471, 0.0365564, 0.1048920, 0.0494506, 0.0918046, 0.1178720, 0.0441359, 0.1363750, 0.0736602, -0.0805816, 0.0205179, -0.0663354, 0.0640431, -0.1153730, -0.0471940, 0.0541421, 0.1932570, -0.0000582, -0.0328812, -0.0047031, -0.0242122, -0.0534006, -0.0183056, 0.0047651, 0.0012003, -0.0000078, -0.0004480, 0.0133289, 0.0094436, 0.0658715, 0.0921485, 0.0982974, 0.1786050, 0.0350417, -0.0549107, 0.1079960, 0.1233640, 0.0770693, 0.0463539, 0.0126832, 0.0454319, 0.0494287, -0.2656240, 0.0429060, -0.0072574, 0.1263380, 0.0647132, 0.0256561, 0.0150112, 0.0622228, 0.0689785, 0.0156020, 0.0018210, -0.0008944, 0.0001501, 0.0082130, 0.0248715, 0.0809315, 0.1128420, 0.1195740, 0.0771873, -0.0253255, -0.0176112, 0.0678290, 0.1804910, 0.0793112, -0.0139162, -0.0187655, -0.1306980, -0.2555850, -0.1015350, 0.0346560, 0.0768857, -0.0798490, -0.1290170, -0.0317353, 0.0099917, 0.1012580, 0.0541224, 0.0047357, 0.0010929, 0.0000379, -0.0006164, 0.0114503, 0.0310040, 0.0542539, 0.0492498, -0.0246844, -0.1965260, 0.0640683, -0.0567091, -0.2072990, 0.0181935, 0.2963190, 0.0765164, -0.0838762, -0.1409750, 0.0689669, -0.0719992, 0.0354339, 0.0240135, 0.0101650, -0.0492408, -0.1981460, -0.1160260, -0.0025589, 0.0119570, -0.0097744, 0.0004457, -0.0002062, -0.0008390, 0.0056326, 0.0054402, 0.1360900, -0.0081055, 0.1075510, 0.0355477, 0.0190435, 0.0996616, 0.1005260, 0.4503200, 0.1892140, -0.2267030, -0.2511090, -0.1029420, 0.2082980, 0.1054450, -0.1976700, -0.2397890, 0.0511864, -0.1934770, -0.2601640, -0.1750610, -0.0650422, 0.0170594, 0.0221937, 0.0044264, 0.0003394, -0.0005412, 0.0027969, 0.0687050, 0.1189550, -0.0960771, -0.0203958, -0.0044994, -0.1144220, 0.1002630, 0.0953772, 0.0058981, -0.0926675, -0.0905359, -0.2134060, -0.0331464, -0.1821950, 0.1279350, -0.2182850, -0.1632590, 0.1007810, -0.1559940, -0.1089140, -0.1073060, 0.0770129, 0.1129780, -0.0014652, 0.0045319, -0.0001813, -0.0017584, 0.0059918, 0.0627310, 0.0612475, -0.0835925, 0.0803345, 0.0017902, -0.0361245, 0.0891506, 0.1621800, 0.0732078, 0.0522748, -0.3945480, -0.2703930, -0.0593118, 0.1073490, 0.3438080, 0.1765550, 0.0841418, 0.3087430, 0.0132303, 0.0955224, 0.1168550, 0.1238010, 0.0103795, -0.0435455, 0.0009208, 0.0001059, 0.0009347, 0.0013549, 0.0243930, 0.0440802, -0.0400066, 0.1055740, -0.0520366, -0.0405021, 0.1005350, 0.0252551, -0.0206683, -0.1420950, -0.5405500, -0.1267040, -0.0400438, 0.0751896, -0.0197668, 0.2210110, 0.0837490, 0.2532850, 0.1344700, 0.0625171, 0.2263180, -0.0522892, -0.0728602, -0.0249496, -0.0020717, 0.0002747, 0.0021245, -0.0013231, 0.0049774, 0.1322820, 0.0104702, 0.0901339, 0.0751718, -0.0140319, -0.0907652, -0.0019077, -0.2279760, -0.2933700, -0.3948210, -0.0549755, -0.1514920, 0.0394531, 0.1043810, 0.0293569, 0.0961295, -0.0545617, 0.1132660, 0.0885303, 0.1647370, -0.0129937, -0.0402915, -0.0475106, -0.0114517, -0.0001516, 0.0045740, 0.0001825, 0.0013440, 0.1463800, 0.0165197, 0.0636088, 0.0594627, 0.0521094, 0.0005693, 0.2094880, -0.1925340, -0.5236160, -0.2354210, -0.2133520, -0.1316140, 0.0335891, 0.1274150, 0.2638800, 0.1188620, 0.2219970, 0.1981740, 0.2628400, 0.2352240, 0.0677164, -0.0740116, -0.0692689, -0.0008750, 0.0002614, 0.0088766, 0.0106986, 0.0020206, 0.1147520, 0.0124749, 0.0919673, 0.1363540, -0.1547920, -0.2009980, 0.2473440, -0.1230200, -0.3591470, -0.3139070, -0.3315250, -0.2003780, -0.1712060, 0.0382259, 0.0406743, 0.1334110, 0.1916220, 0.2558270, 0.1513380, 0.0568185, -0.0012608, -0.1262590, -0.1082790, -0.0233468, 0.0004009, 0.0036164, 0.0326058, 0.0380373, -0.0888649, -0.0081448, 0.0160579, 0.1993170, 0.0744097, 0.3162800, 0.1999160, 0.1638260, -0.1633560, -0.2769070, -0.2662230, -0.1566650, -0.2873210, -0.2068360, 0.1182860, 0.1789890, 0.1576390, 0.1732180, 0.1164520, 0.0098314, 0.0855132, -0.1849120, -0.1594330, -0.0486905, 0.0002076, 0.0014728, 0.0466489, 0.0586801, -0.1717250, -0.0697232, 0.0872190, 0.1929470, 0.2316550, 0.0980050, 0.2343550, 0.0316372, -0.0722735, -0.2112250, -0.1738810, -0.2613420, -0.1535850, 0.1909430, 0.2904210, 0.2380540, 0.0336489, 0.0380882, 0.0837708, 0.0214295, -0.0051036, -0.2330900, -0.0663136, -0.0177545, 0.0002987, -0.0001849, 0.0230597, 0.0714400, -0.0794954, -0.0339958, 0.0105479, 0.1533090, 0.0269784, 0.0795502, 0.2660020, 0.2526500, -0.0273896, -0.3296120, -0.4087940, -0.3715860, -0.0115566, 0.3730050, 0.3121010, 0.4947610, 0.2800000, 0.1064550, 0.1102270, -0.0287410, -0.0944457, -0.1598100, -0.0215123, -0.0113899, -0.0003631, 0.0004253, 0.0013448, 0.0295699, -0.0018796, 0.0807820, -0.0795103, 0.0598487, 0.1395450, 0.0768864, 0.0970074, 0.2685800, 0.0873447, -0.3788620, -0.4207940, -0.2325270, 0.3445380, 0.3337710, 0.3546570, 0.2869250, 0.0527314, 0.0946565, 0.1254440, -0.1054140, -0.0196651, -0.0991317, -0.0467896, -0.0015962, 0.0003692, 0.0004882, -0.0189378, -0.0982134, -0.0481701, -0.0090746, -0.1051640, -0.1261630, 0.0329301, 0.1016570, -0.1911300, -0.2204640, -0.3086190, -0.3565340, -0.1124620, 0.0479478, 0.4934550, 0.2952700, 0.2092930, 0.2187990, 0.0020293, -0.0520794, -0.0112000, -0.0621022, 0.0374708, 0.0636739, -0.0167237, -0.0001756, -0.0005421, -0.0005433, -0.0684254, -0.1519000, -0.0917277, -0.0727298, -0.1092220, -0.1559330, -0.0115914, -0.2321140, -0.2732110, -0.0641454, -0.1669420, -0.3104470, -0.1373810, 0.3664580, 0.5863480, 0.0773042, 0.0326565, 0.1432420, 0.1512180, -0.0282117, 0.0185793, -0.0571064, 0.1249260, 0.0912161, -0.0015258, 0.0005570, -0.0001559, 0.0004298, -0.0713065, -0.0897716, -0.1067030, -0.1046860, -0.2933850, -0.2411940, -0.2787610, -0.3719840, -0.4095110, -0.2821010, -0.1380090, -0.1140960, 0.0409303, 0.3077410, 0.4688610, 0.1265170, 0.1124780, -0.0577327, 0.0482873, -0.0753602, -0.0905039, 0.0339745, 0.1004420, 0.0974285, 0.0115226, -0.0000559, -0.0001854, -0.0001321, 0.0013794, 0.0060547, -0.0172547, 0.0091940, -0.0347595, -0.1413410, -0.1597320, -0.3296710, -0.0848181, 0.0743231, -0.1402700, 0.0655312, 0.4720970, 0.3089690, 0.2800160, 0.2857510, 0.1523340, 0.0251301, 0.1534370, 0.0667996, 0.0192715, 0.1225200, 0.0949883, 0.0576700, 0.0058263, 0.0001156, -0.0000683, -0.0001557, 0.0033708, 0.0067842, 0.0062852, 0.0250286, 0.0351408, 0.0536964, -0.0704456, -0.0124955, 0.2158700, 0.1549110, -0.0043537, 0.1917500, 0.2578940, 0.2109980, 0.3189560, 0.4535440, 0.1440590, -0.0180222, 0.1386580, 0.0565116, 0.1058940, 0.1353610, 0.0089728, -0.0258493, -0.0066673, 0.0000068, 0.0007617, -0.0003092, 0.0008389, -0.0004800, -0.0034686, -0.0028186, 0.0169235, 0.0363708, 0.0383238, 0.0329718, 0.0944943, 0.1293660, 0.0421673, 0.1230220, 0.1673420, 0.1428800, 0.2056070, 0.1926120, 0.2156330, 0.2891210, 0.1743600, 0.1570300, 0.1208240, 0.0835783, 0.0402637, -0.0054371, -0.0072814, -0.0002318, 0.0000867, 0.0001786, -0.0002199, 0.0008592, 0.0016225, 0.0220818, 0.0220685, 0.0037727, 0.0025773, 0.0395120, 0.0111333, 0.0360302, 0.0179314, -0.0041078, 0.1526410, 0.2222090, 0.2137500, 0.1650070, 0.1090390, 0.0707608, 0.1056080, 0.0866247, 0.0268154, 0.0039133, 0.0002306, -0.0001254, -0.0000080, 0.0003831, -0.0001001, -0.0001783, 0.0001863, 0.0001246, -0.0000340, 0.0001213, 0.0009966, 0.0097768, 0.0083832, -0.0035286, -0.0150501, -0.0186858, -0.0181289, -0.0221998, 0.0075657, 0.0219942, 0.0057326, -0.0023483, 0.0128417, 0.0087944, 0.0164822, 0.0045891, 0.0052193, 0.0000926, 0.0002130, -0.0001960, 0.0005525, 0.0001398, -0.0000272, -0.0002554, 0.0005508, 0.0000284, -0.0004033, 0.0000384, 0.0000184, -0.0001206, 0.0004599, 0.0005961, 0.0002611, 0.0000199, 0.0000600, -0.0004450, 0.0002207, 0.0001837, 0.0000664, -0.0000227, 0.0000359, 0.0007064, -0.0000875, -0.0007018, 0.0001891, 0.0000205, -0.0003368, -0.0004675, -0.0003718, 0.0001709, 0.0006115, -0.0000638, -0.0004723, 0.0003192, 0.0001533, -0.0003235, 0.0000260, 0.0002145, 0.0012081, -0.0004845, -0.0009765, -0.0001547, 0.0012262, -0.0004298, -0.0197973, -0.0376382, -0.0055759, -0.0011590, -0.0006007, -0.0007037, -0.0010245, -0.0004516, 0.0027224, 0.0040432, 0.0003774, 0.0003240, -0.0004409, -0.0005986, -0.0003334, -0.0005312, 0.0001020, 0.0000327, 0.0000078, -0.0001883, 0.0003152, 0.0022878, 0.0129078, 0.0378763, 0.0459490, 0.0525752, 0.0078062, -0.0492752, 0.0057932, -0.0812424, -0.0594270, 0.0003128, -0.0335422, -0.0420135, -0.0116664, 0.0024013, 0.0010212, 0.0028557, 0.0002641, -0.0002948, -0.0006798, -0.0005485, -0.0003690, 0.0000615, -0.0051529, -0.0013732, 0.0019583, -0.0309693, -0.0337103, -0.0491810, -0.0399045, 0.0171253, -0.0074354, 0.1174570, -0.0263261, -0.0985831, 0.0198049, 0.0950364, 0.0833939, -0.0427086, -0.1415570, 0.0052392, -0.0174229, 0.0481859, 0.0039867, -0.0050296, 0.0287101, -0.0167173, 0.0071838, 0.0001482, 0.0001604, -0.0000313, -0.0169403, -0.0071824, -0.0017334, -0.0185041, 0.0155941, 0.0418952, 0.0331395, 0.1134460, 0.1567690, 0.0875843, 0.0777503, -0.0282624, -0.0717069, -0.1968780, -0.1216710, -0.2209710, -0.3027090, 0.0304500, 0.0516297, 0.0398568, -0.0179948, 0.0135150, 0.0134382, -0.0167356, -0.0133927, 0.0100550, 0.0000789, -0.0003594, -0.0024343, -0.0072016, 0.0289248, -0.0397472, -0.0133769, 0.0026748, -0.0050415, 0.0111137, 0.1293660, 0.0027575, -0.0316801, -0.0488066, 0.2458010, 0.0160933, -0.0645984, -0.1779310, 0.0314175, 0.1083280, 0.0683436, 0.0111393, -0.0375746, 0.0782137, 0.0299587, -0.0422406, 0.0313277, 0.0183868, -0.0004876, -0.0002943, -0.0079663, 0.0208283, 0.0615056, -0.0326623, -0.0752200, -0.1790190, -0.1375830, -0.1733700, -0.3655360, -0.2044530, -0.1423720, -0.1614690, -0.1002480, -0.0521678, 0.0174866, -0.1537970, -0.3095290, -0.3976520, -0.3168230, -0.2294250, -0.1539640, -0.0368438, -0.0222666, -0.0408349, -0.0046592, 0.0063456, 0.0000815, 0.0008570, 0.0011176, 0.0137028, 0.0382508, -0.1083540, -0.0892895, -0.1227590, -0.1049950, -0.2717580, -0.4951960, -0.2251090, -0.2264790, -0.2035860, -0.1034660, -0.2583160, -0.0677373, -0.1219760, -0.4381100, -0.6054230, -0.3358850, -0.2022910, -0.0323498, -0.1386180, -0.0131822, 0.0195379, 0.0440035, 0.0040594, 0.0026334, 0.0015101, -0.0042509, -0.0184746, -0.0168431, 0.0101372, -0.0096136, -0.1415010, -0.1728290, -0.0319800, -0.1706440, -0.2290210, -0.2443230, 0.0062226, -0.1199430, -0.0281813, -0.0916402, -0.0815611, -0.3941970, -0.1301240, -0.1327350, -0.1950600, -0.0907795, -0.0116969, 0.0463184, 0.1125280, -0.0283643, -0.0062710, -0.0001533, -0.0003957, -0.0081192, -0.0302665, -0.0897833, 0.0027961, -0.2423060, -0.1811440, -0.3484520, -0.2875040, -0.2108220, -0.2810580, -0.0726798, -0.0908849, -0.3061330, -0.2596330, -0.0410547, -0.1439400, -0.1997390, -0.1033320, 0.0688754, -0.0548462, -0.0488244, -0.0554746, 0.0579923, -0.0239759, -0.0304855, -0.0017331, -0.0005603, 0.0003197, -0.0163220, -0.0173487, -0.0970536, 0.0091702, -0.2335670, -0.1147840, -0.2739560, -0.1377530, -0.2737320, -0.1637100, -0.1070890, -0.1351390, -0.2260330, -0.1447390, -0.0377265, 0.0104403, -0.0618823, -0.0527852, -0.0167974, 0.0271504, -0.0151659, -0.1986240, 0.0536242, -0.0119057, -0.0018885, -0.0059186, -0.0002317, 0.0012446, -0.0085639, -0.0189351, -0.2031430, -0.0791985, -0.0264828, -0.1412650, -0.0979155, -0.2530410, -0.1707960, -0.2400200, -0.1760520, -0.2218100, -0.2250180, -0.3302140, 0.1901250, -0.1294730, -0.1155610, 0.1691120, -0.0583444, 0.0462064, -0.1144000, -0.2391120, -0.1155920, 0.0066690, -0.0430444, -0.0061735, -0.0004231, -0.0001968, -0.0040942, -0.0474633, -0.2677380, -0.1882110, -0.1592150, -0.0673405, 0.0951482, -0.0833222, 0.0456509, 0.0894015, -0.0491191, -0.0983792, -0.3403760, -0.4040220, 0.0401053, -0.3012050, -0.2545210, -0.2217720, -0.1646560, -0.1615670, 0.0274189, -0.3188490, -0.0563606, 0.0119026, -0.0616271, -0.0050084, -0.0002787, -0.0004310, -0.0027190, -0.0540183, -0.3255170, -0.0708266, 0.0700126, -0.0018811, 0.1056000, -0.0608881, 0.2235890, 0.0963179, 0.1646730, 0.0079036, -0.2909840, -0.2008500, -0.0831406, -0.2439740, -0.2287980, -0.2623740, -0.2843340, -0.0650830, 0.0220978, 0.1343990, 0.1481740, 0.0232990, -0.0092185, 0.0082894, 0.0003737, -0.0012942, -0.0011405, 0.0035286, -0.1305780, 0.1220630, 0.2793250, 0.2766080, 0.1283410, 0.2789990, 0.1553070, 0.2467160, 0.3582700, 0.0439109, -0.1857700, -0.2231080, 0.1132170, -0.0572236, -0.2103160, -0.2458500, -0.2300370, -0.0046026, 0.2682450, 0.1607920, 0.1939090, 0.0762600, 0.0281807, 0.0007632, 0.0002366, -0.0005412, 0.0053114, 0.0905809, 0.0669078, 0.2672550, 0.2561670, 0.1431550, 0.1854240, 0.4037790, 0.4050240, 0.3421050, 0.3039940, 0.1927580, 0.0863691, -0.0182177, 0.0945309, 0.2524190, -0.2102570, -0.0459786, -0.0676628, 0.0468042, 0.1094220, 0.0739690, 0.1570770, 0.1386130, 0.0564417, 0.0117999, -0.0002783, -0.0004907, -0.0027242, 0.0897392, 0.0797557, 0.2151510, 0.2299890, 0.3184200, 0.2238410, 0.2145920, 0.3357800, 0.4149290, 0.2395140, 0.0349503, 0.0502357, 0.3427030, 0.3870590, 0.4083040, 0.2099160, 0.1318990, 0.1933050, 0.2846820, 0.0669926, 0.1420840, 0.1428450, 0.1754310, 0.0714201, 0.0227779, 0.0004892, -0.0002768, 0.0135212, -0.0018478, 0.0966271, 0.3375360, 0.2528910, 0.1442870, 0.1205800, 0.1272970, 0.2378360, 0.3282220, 0.0350198, 0.0038352, 0.2050340, 0.2306090, 0.2633890, 0.1599710, 0.4582270, 0.1203870, 0.1489770, 0.1647090, 0.1362260, 0.0707323, 0.0220173, 0.1251580, 0.0015385, 0.0151191, -0.0015741, -0.0001428, 0.0061939, -0.0207509, 0.1598330, 0.1836900, 0.2219540, 0.1878010, 0.1752350, 0.1125430, 0.1393880, 0.1232190, 0.2480190, 0.2036680, 0.2805570, 0.1279230, 0.4047900, 0.2973190, 0.3394710, 0.1298590, 0.0243133, 0.1529680, 0.0313921, 0.2000620, 0.1125490, 0.0928660, -0.0094717, 0.0098877, -0.0000341, -0.0033369, -0.0031525, -0.0286355, 0.1019320, 0.0389964, -0.0518536, 0.1629610, 0.0140847, 0.0235198, 0.1819380, 0.2336360, 0.0679406, 0.0545031, 0.2270480, 0.2656600, 0.2142810, 0.3310400, 0.2767590, -0.0436694, 0.1058980, 0.1205630, 0.0215201, 0.0538848, 0.0322080, 0.0833341, 0.0206040, 0.0008258, -0.0001322, -0.0043882, -0.0000077, 0.0603565, 0.0442898, -0.0498190, -0.2341500, 0.1064230, 0.0532332, 0.1087910, 0.0972632, 0.1147730, 0.0657259, -0.1701490, -0.0706886, 0.0805733, 0.0425720, 0.0531803, 0.1146730, 0.0723222, 0.2178870, 0.2624850, 0.0112133, 0.0081321, 0.0264654, 0.0281278, 0.0123066, -0.0003248, -0.0000805, 0.0007279, 0.0031602, 0.0839224, 0.0752357, 0.0141155, -0.1225040, -0.0720064, -0.0759666, 0.0101301, -0.1153300, -0.1217430, -0.0039613, -0.1290080, -0.0596971, -0.0402155, -0.0995366, 0.0480745, 0.0601125, 0.1617130, 0.2038070, 0.1003820, 0.0810857, 0.0838161, -0.0344226, 0.0293826, 0.0065212, 0.0000928, -0.0000570, 0.0000568, 0.0041912, 0.0524475, -0.0211094, -0.0275318, -0.0843559, 0.0037299, -0.0908244, -0.0642875, 0.1210680, 0.1583420, 0.2162460, 0.0187883, -0.0760248, 0.0578317, -0.0228876, -0.1637010, -0.0703283, 0.1077680, 0.0903903, 0.2262320, -0.0354680, -0.0931918, -0.0524544, -0.0339206, 0.0030859, 0.0001722, 0.0000637, -0.0001695, 0.0013376, -0.0024891, -0.0295475, -0.0852586, -0.0910377, -0.0483219, -0.0925923, -0.1222290, -0.0942003, 0.0310571, -0.0406281, -0.2515550, -0.1923650, -0.2618880, -0.3474130, -0.4804810, -0.1922130, -0.1739640, -0.0875716, 0.0266354, -0.1610960, -0.1816300, -0.1049440, -0.0085288, 0.0024784, -0.0002708, 0.0001292, 0.0001575, -0.0003607, -0.0303793, -0.0458210, -0.0733950, -0.1218950, -0.0817467, -0.1884940, -0.1993340, -0.2482410, -0.1644770, -0.3356560, -0.2530410, -0.3433290, -0.1550340, -0.1450440, -0.2753160, -0.2108430, -0.2695760, -0.2012380, -0.1473620, -0.1680360, -0.1692400, -0.0426750, 0.0043059, 0.0031802, 0.0001790, -0.0000928, -0.0003616, -0.0001711, -0.0002009, -0.0044921, -0.0481050, -0.0724026, -0.0699598, -0.1752600, -0.2884230, -0.2148820, -0.1255630, -0.2775710, -0.3084540, -0.3143140, -0.1845630, -0.1807730, -0.3082140, -0.4136490, -0.4246680, -0.2066760, -0.1383570, -0.0725443, -0.0514575, -0.0239186, 0.0024743, 0.0023078, -0.0005125, -0.0009023, -0.0002875, 0.0000140, 0.0001492, -0.0013156, -0.0409727, -0.0677514, -0.0718878, -0.0811619, -0.0762396, -0.0781162, -0.1201030, -0.1204550, -0.1065470, -0.1489010, -0.1334820, -0.1028560, -0.0487357, -0.1177580, -0.1155790, -0.0954975, -0.0688886, -0.0356968, -0.0048368, -0.0028249, -0.0000872, 0.0001361, 0.0000317, -0.0005373, 0.0001808, -0.0002091, -0.0000173, 0.0000700, 0.0001435, -0.0050708, -0.0295601, -0.0266619, -0.0055428, -0.0108072, -0.0079372, -0.0073681, -0.0089195, -0.0307361, -0.0072873, -0.0059969, -0.0113306, -0.0364477, -0.0128647, -0.0043673, -0.0233898, -0.0318604, -0.0044236, -0.0000991, -0.0005359, 0.0001103, 0.0000362, 0.0000942, 0.0003579, -0.0005421, 0.0006940, -0.0004797, -0.0004616, -0.0000782, 0.0003382, -0.0004583, -0.0000085, 0.0000507, 0.0005370, 0.0002323, -0.0002062, -0.0000222, 0.0001004, -0.0004463, 0.0003327, -0.0003745, 0.0000168, -0.0002046, 0.0006745, -0.0009021, 0.0004269, -0.0001008, 0.0001605, -0.0011007, 0.0003919, -0.0002473, 0.0002759, -0.0007279, 0.0004937, -0.0004388, -0.0005034, -0.0056848, -0.0109616, -0.0278574, -0.0127563, -0.0191908, -0.0139841, -0.0154768, -0.0165792, -0.0125303, -0.0024029, -0.0018868, -0.0011925, -0.0000810, -0.0003350, -0.0003496, -0.0005168, -0.0046945, -0.0064580, -0.0001795, -0.0001444, -0.0000274, 0.0002743, -0.0002029, -0.0003609, -0.0001858, 0.0000980, -0.0001949, -0.0003261, -0.0052721, -0.0224218, -0.0458829, -0.0569066, -0.0887961, -0.0886830, -0.1050070, -0.0868412, -0.0478937, -0.0232201, -0.0086473, 0.0002751, -0.0018368, 0.0006099, -0.0014858, -0.0041433, -0.0063055, -0.0055444, -0.0011381, 0.0002197, 0.0002551, 0.0002038, -0.0002291, 0.0000783, 0.0007619, 0.0002197, 0.0008609, -0.0064093, -0.0299814, -0.0284369, -0.0823399, -0.0977628, -0.0757927, -0.1724160, -0.1771690, -0.1086230, -0.0475259, -0.0161774, -0.0042954, 0.1336580, 0.1718500, 0.1372300, 0.0939698, 0.0330596, -0.0020111, -0.0070748, 0.0028372, 0.0002824, 0.0000295, 0.0005321, 0.0003205, -0.0000714, -0.0005702, -0.0003148, -0.0058558, -0.0258703, -0.0559794, -0.0363730, -0.0561776, -0.0108533, 0.0135681, 0.0171350, -0.0215831, -0.0613324, -0.1066730, 0.0320843, 0.1429100, 0.1312290, 0.1041450, 0.1358630, 0.1401690, 0.1863780, 0.1438290, 0.0927124, 0.0511920, 0.0238870, 0.0062490, -0.0012834, -0.0000665, 0.0004233, -0.0009874, -0.0085266, -0.0557711, -0.0332323, -0.0532971, 0.0770083, 0.1745400, 0.2993370, 0.2104650, -0.0643290, -0.2462470, -0.5322100, -0.3071670, -0.2342000, 0.0299961, 0.1141540, 0.1406290, 0.0226749, 0.0758927, 0.1224040, 0.1357890, 0.1028920, 0.0792542, 0.0448418, 0.0032710, 0.0035808, -0.0003334, 0.0000402, -0.0028737, -0.0165531, -0.0593169, 0.0538252, 0.1232120, 0.0658446, 0.1724350, 0.2229540, 0.0820864, -0.0859979, -0.4069780, -0.8176590, -0.5252360, -0.0561583, 0.0593811, 0.0383479, 0.1516450, 0.1170820, 0.0269345, 0.0847967, 0.1058880, 0.1161600, 0.0952510, 0.0537468, 0.0320012, 0.0096436, 0.0003825, 0.0006207, -0.0013645, -0.0187770, -0.0649375, 0.0865766, 0.1840270, 0.2217900, 0.1574430, 0.1902750, 0.1768430, 0.1185210, -0.3261240, -0.9091770, -0.5028530, 0.0080976, 0.3030100, 0.1534890, 0.0673144, 0.0764839, -0.0595858, -0.1338390, 0.0483789, 0.1424480, 0.0992691, 0.0430419, 0.0339603, 0.0010404, -0.0001396, 0.0068686, 0.0064207, -0.0028550, -0.0184596, 0.1443570, 0.0916766, 0.0703412, -0.0130003, 0.2300510, 0.2908760, 0.1843790, -0.4368850, -0.6451370, -0.3370690, 0.0615341, 0.1947130, 0.1884000, -0.0603574, -0.1896460, 0.1354610, -0.0099074, -0.0225054, 0.1919230, 0.1255640, 0.0734596, 0.0024807, -0.0048288, 0.0004167, 0.0104540, 0.0219289, -0.0045252, 0.0241604, 0.0273870, 0.0945053, -0.0467251, 0.1464610, 0.2240630, 0.4845980, 0.2566570, -0.3717230, -0.7749680, -0.2926870, 0.0545738, 0.2375070, -0.1248900, -0.1798540, -0.2761530, 0.0468929, -0.0018989, -0.1477490, 0.0810112, 0.0602410, 0.0737234, 0.0174486, 0.0025535, -0.0000075, 0.0103596, 0.0279821, 0.0037175, 0.0101244, 0.0318628, -0.0083246, -0.0139244, 0.1213150, 0.3650410, 0.6245640, 0.4694080, -0.1463310, -0.6357210, -0.5334020, 0.0086644, 0.0057432, -0.2098040, -0.2343560, -0.0973127, -0.1235470, -0.0663639, -0.1391020, -0.1740590, -0.0016282, 0.0975639, 0.0185902, 0.0016636, 0.0006387, 0.0081683, 0.0615535, 0.0581752, 0.0188124, 0.1470380, 0.1950560, -0.0534705, -0.0433208, 0.2759180, 0.5299420, 0.5908180, -0.1581940, -0.6877680, -0.3689120, -0.0815175, 0.0902793, -0.1400590, -0.0638222, -0.1512630, -0.2518040, -0.1173770, -0.1821260, -0.0402193, -0.0081930, 0.0266497, 0.0130713, 0.0006649, 0.0004006, 0.0028833, 0.0513305, 0.0667085, 0.0244368, 0.0934654, 0.0897559, 0.1950850, 0.1130810, 0.3055950, 0.4403620, 0.4111520, -0.1222860, -0.3835030, -0.4430160, 0.1973120, 0.1252280, -0.1039580, -0.0547352, 0.0858757, 0.2107080, -0.0147975, 0.0383955, -0.0804669, -0.1386020, -0.0021315, 0.0263760, 0.0020529, 0.0002501, 0.0015504, 0.0353598, 0.0235834, 0.0966568, 0.2417990, 0.1032390, 0.1590290, 0.1701530, 0.1477790, 0.1846310, 0.1706470, -0.0915340, -0.1831660, -0.2479110, -0.1073370, -0.3473790, -0.1955870, -0.0497343, -0.0600425, 0.2125130, 0.1029430, 0.0591140, -0.1076990, -0.0388456, -0.0246712, -0.0065673, -0.0033114, 0.0013277, 0.0003227, 0.0277871, -0.0112543, 0.0612845, 0.2662890, 0.1839180, 0.1340940, 0.3163000, 0.3325130, 0.0106062, -0.0819405, -0.1096510, -0.1754590, -0.1209360, -0.0298844, -0.1190820, -0.0616378, -0.0475344, 0.0768368, -0.0369066, -0.0197311, 0.0404482, 0.0357344, 0.0670623, -0.0624482, -0.0085829, 0.0000414, -0.0001977, -0.0001448, 0.0123863, 0.0310544, 0.0719519, 0.0531991, 0.1818160, 0.1563970, 0.2001530, 0.1440020, 0.0500580, 0.0076485, -0.0825377, -0.0767042, -0.0976028, 0.0274361, -0.1942740, -0.1546550, -0.0096191, 0.1150170, -0.1783360, -0.1280070, -0.0333366, 0.0213245, -0.0105110, -0.0382126, 0.0294582, -0.0004545, -0.0008241, -0.0000443, -0.0018341, 0.0501952, 0.0131629, -0.0767161, 0.0372048, -0.0479574, 0.1257680, 0.0539687, -0.1418020, -0.3007010, -0.1196570, -0.2788400, -0.0433113, 0.0745736, -0.0098299, -0.2606170, -0.2814590, 0.1104890, 0.1186330, 0.0803106, -0.0542568, -0.0109646, 0.0096588, 0.0281236, 0.0207174, 0.0002063, 0.0002917, 0.0005931, 0.0182389, 0.0170142, 0.0455665, 0.0173789, -0.0703060, -0.1042440, -0.1168220, -0.0619326, -0.1870110, -0.2699660, -0.2299990, -0.2880170, -0.1536940, -0.2201600, -0.0449494, -0.1960610, -0.0122398, 0.0176845, 0.0918352, -0.0559870, -0.1158050, -0.0245408, 0.0192719, 0.0348811, 0.0103977, -0.0003962, -0.0000491, -0.0006594, 0.0098856, -0.0120906, 0.0402239, 0.0312602, -0.2359410, -0.3158910, -0.2163730, -0.0949237, -0.0561441, -0.1229890, -0.2498550, -0.2425630, -0.0361194, -0.2128990, -0.1537790, -0.1759420, -0.0781216, -0.0709198, -0.0711236, -0.0878725, -0.1839450, -0.0650578, 0.0358899, 0.0072472, 0.0002914, -0.0002155, 0.0002622, 0.0003444, -0.0035530, -0.0477775, -0.0396409, -0.0539125, -0.1276010, -0.1586000, -0.1025850, -0.1383990, -0.1521360, -0.1111860, -0.2487890, -0.1233180, -0.0581852, -0.1783010, -0.3060250, -0.1199770, -0.0854055, -0.0593689, 0.0108675, -0.0054929, -0.1496120, -0.0469091, 0.0261497, 0.0253767, 0.0000093, 0.0004178, 0.0005973, 0.0003710, -0.0040600, -0.0511514, -0.0948191, -0.1287830, -0.0745654, -0.0758340, 0.0323261, -0.0960140, -0.1533140, -0.1819640, -0.0908638, 0.0304448, -0.1462390, 0.0456313, -0.1518940, 0.0537853, 0.1150860, 0.0456467, 0.0100739, -0.0195431, 0.0415407, -0.0027392, -0.0630423, -0.0153011, 0.0003388, -0.0007876, -0.0000992, 0.0001657, -0.0032268, -0.0401089, -0.0488190, -0.1143890, -0.0895820, -0.0758616, 0.0052372, -0.1332290, -0.1418410, -0.0652802, -0.2025980, -0.1172180, 0.0563454, 0.0156528, 0.0187078, 0.0925147, 0.1674760, 0.0448318, 0.1149860, 0.1669950, 0.0182037, 0.0304103, 0.0091812, 0.0327882, 0.0004342, -0.0002649, 0.0001612, 0.0000797, -0.0020857, -0.0188572, -0.0271945, -0.0293655, -0.0450038, -0.0528624, 0.0086007, -0.1367510, -0.2588310, -0.2715950, -0.2745120, 0.0544152, 0.3244100, 0.1561700, -0.0326601, 0.1061300, 0.1407730, 0.0682678, 0.0913622, 0.1749470, -0.0403085, -0.0023450, 0.0202758, 0.0210171, 0.0094875, -0.0000114, -0.0004674, 0.0005932, -0.0016145, -0.0024407, 0.0083153, 0.0123600, 0.0015724, -0.0155338, -0.0439018, -0.0029590, 0.0299612, -0.1236620, 0.0542068, 0.0605552, 0.2662520, 0.1134930, 0.2069910, 0.0914320, 0.0290190, -0.0815314, 0.0283727, 0.0692369, -0.1466870, -0.1008990, -0.0638760, 0.0250111, 0.0079409, -0.0003426, 0.0001553, -0.0007887, -0.0020706, -0.0029888, -0.0005413, 0.0033577, 0.0022031, 0.0502812, -0.0057455, -0.0812786, -0.1190500, -0.0123928, 0.1263200, 0.1939390, 0.1893380, 0.1162750, -0.0223037, 0.2129750, 0.0892918, -0.0090753, -0.0494365, -0.0814096, -0.1242120, -0.1325160, -0.0326112, -0.0003698, 0.0005024, 0.0000514, -0.0000350, 0.0007642, -0.0004922, 0.0013114, 0.0067760, -0.0328403, -0.0630177, -0.0569549, -0.0499326, -0.1809750, -0.1632850, -0.0281987, -0.0442305, 0.0021436, 0.0227658, 0.1750860, 0.1122370, 0.2037500, 0.1276600, -0.0455841, -0.0832545, -0.0645075, 0.0068830, -0.0149654, -0.0058162, -0.0002977, -0.0001077, 0.0000419, 0.0000282, 0.0000469, 0.0000266, -0.0001363, -0.0020732, -0.0397776, -0.0549250, -0.0474535, -0.0101898, -0.0394490, -0.0955428, -0.0540722, -0.0750306, -0.1031620, -0.1563730, -0.0003266, -0.0963053, -0.1345400, -0.1686650, -0.0419562, -0.0802511, -0.0774474, -0.0121834, -0.0174844, -0.0046847, -0.0001030, 0.0001629, 0.0004579, -0.0000296, 0.0003363, 0.0003556, 0.0007938, -0.0001504, 0.0000444, -0.0007855, -0.0085856, -0.0072826, 0.0040406, 0.0128958, 0.0060018, 0.0048643, 0.0180235, -0.0416102, -0.0509749, -0.0063403, -0.0018681, -0.0429016, -0.0166033, 0.0054553, -0.0016305, 0.0057409, 0.0047315, 0.0005921, -0.0002622, -0.0000347, -0.0001571, -0.0007030, 0.0000063, 0.0001432, -0.0000038, -0.0003072, -0.0001021, 0.0001514, 0.0001889, -0.0003917, -0.0001433, 0.0004712, -0.0000621, 0.0002919, 0.0002831, -0.0004494, 0.0001229, 0.0008700, -0.0001847, -0.0002389, -0.0000034, -0.0001851, 0.0000672, 0.0003241, -0.0004824, -0.0000632, -0.0002355, -0.0005135, -0.0000029, -0.0007277, 0.0002739, 0.0001793, 0.0001577, 0.0003237, -0.0003955, -0.0004523, -0.0013957, -0.0023609, -0.0031237, -0.0104967, -0.0108342, -0.0107835, -0.0016438, 0.0077007, -0.0050285, 0.0108862, -0.0036789, -0.0081749, -0.0151869, -0.0188739, -0.0114226, -0.0024255, 0.0001152, -0.0000737, 0.0004986, 0.0003167, -0.0005235, 0.0003471, -0.0003053, -0.0005395, 0.0001512, -0.0004621, -0.0008382, -0.0061490, -0.0099753, -0.0308795, -0.0432497, -0.0414443, -0.0383061, -0.0034575, 0.0444406, 0.0000276, -0.0391118, -0.0375874, -0.0401626, -0.0869260, -0.0889804, -0.0729588, -0.0619101, -0.0406623, -0.0185219, -0.0067895, 0.0000197, -0.0003167, 0.0001545, -0.0001621, 0.0001946, -0.0000455, -0.0011001, -0.0083976, -0.0096344, -0.0343839, -0.0486756, -0.0663864, -0.1065110, -0.0817624, -0.0933680, -0.0308180, 0.0401855, 0.1553580, 0.0606375, 0.0817035, 0.0535376, -0.0296235, -0.0358813, -0.0408549, -0.0626277, -0.0604124, -0.0764963, -0.0372935, 0.0086914, 0.0031538, -0.0003505, -0.0004166, 0.0002469, 0.0005123, 0.0004650, -0.0143675, -0.0132413, -0.0285369, -0.0137404, -0.0244763, 0.0291260, 0.0169379, 0.0821945, 0.1822640, 0.2867130, 0.2260720, 0.1407280, 0.1458350, 0.1820990, 0.1103740, -0.0227853, -0.0324837, -0.0600725, 0.0164379, -0.0516143, -0.0446078, -0.0039682, -0.0018538, -0.0058122, 0.0001222, 0.0003725, -0.0005857, 0.0013516, -0.0551853, -0.0790231, -0.1056380, -0.1278010, -0.0845403, -0.0692946, -0.0323515, 0.0258807, -0.0211289, 0.0791189, 0.0336691, 0.1497290, 0.2662930, 0.1339850, 0.1890430, 0.0750216, -0.0092874, 0.2022760, 0.1522620, 0.0414434, -0.0421887, -0.0468223, -0.0185166, -0.0148931, 0.0002991, 0.0003189, -0.0025403, -0.0058930, -0.0841457, -0.1042080, -0.1020430, -0.2021870, -0.2106160, -0.1770760, -0.1358500, -0.1817990, -0.1262930, -0.0563800, 0.2273500, 0.1361890, 0.1860110, 0.1581630, 0.4157800, 0.1246150, 0.0656634, 0.2511570, 0.1024790, -0.0616987, -0.1251710, -0.0763128, -0.0228941, -0.0166082, 0.0003287, 0.0008127, 0.0005573, -0.0109915, -0.0722399, -0.0811807, -0.0926916, -0.1517870, -0.1380940, -0.2091890, -0.1284530, -0.2036250, -0.1203040, -0.2102710, 0.1086170, 0.1166450, 0.2791180, 0.2606820, 0.1769050, 0.3223850, 0.0958275, 0.1249460, 0.0742300, -0.0332797, -0.1585950, -0.0556583, -0.0223442, -0.0030887, 0.0007945, 0.0001379, -0.0035095, -0.0284003, -0.0381452, -0.1373880, -0.1494160, -0.1996140, -0.2159730, -0.2406800, -0.3247020, -0.1495750, 0.0417056, -0.2863460, 0.0457234, 0.0950083, 0.4177240, 0.2708410, 0.1160350, 0.0949681, 0.2050940, 0.0228491, 0.1225060, -0.0947314, -0.1789590, -0.0810661, -0.0161896, -0.0016573, 0.0001089, -0.0004162, -0.0057266, -0.0231137, -0.0610402, -0.0895059, -0.2074650, -0.2559430, -0.2391450, -0.0397126, -0.0444899, -0.1512770, -0.0568738, -0.1727590, -0.1834880, -0.1043830, 0.3163110, 0.3721770, 0.3688450, 0.2620990, 0.1730380, -0.0323673, 0.0621488, -0.0463638, -0.1495870, -0.0946252, -0.0503908, 0.0001779, -0.0004346, -0.0026796, -0.0100559, -0.0110925, -0.1312810, -0.1083260, -0.0352747, -0.2429350, -0.0677984, -0.0124996, -0.1611990, -0.1454580, -0.1815090, -0.2518790, -0.3201320, -0.1313820, 0.1758730, 0.5904990, 0.5265800, 0.1820470, -0.0563652, 0.0868185, 0.1415620, -0.1412040, -0.1573660, -0.0429683, -0.0217214, 0.0003653, -0.0000347, 0.0016507, -0.0071712, -0.0412793, -0.0910917, -0.0997902, 0.1813620, -0.1661020, -0.0032148, -0.0651782, -0.0721636, 0.0239397, 0.0557743, -0.0505954, -0.4574210, -0.3893840, -0.1550300, 0.3297000, 0.4564350, 0.3842910, 0.0907111, 0.0481423, -0.0474566, -0.0887546, -0.1098170, -0.0334726, -0.0033945, -0.0001342, -0.0000320, -0.0015789, -0.0033445, -0.0499989, 0.0401256, -0.0121071, 0.1537360, -0.0360977, 0.0623163, 0.0496778, 0.0129278, -0.1206340, 0.0066639, -0.2685740, -0.5164230, -0.4094930, -0.2589050, -0.1136660, 0.1034820, 0.2517560, 0.1866910, -0.0345372, -0.0487331, -0.1595730, -0.1791820, -0.0626878, -0.0093584, 0.0006057, 0.0004310, -0.0001747, -0.0028504, -0.0326875, 0.1065180, 0.1208520, 0.0891039, 0.0593346, -0.0146744, -0.2382530, -0.1090610, -0.2541330, -0.1309420, -0.3982500, -0.3443460, -0.3338620, -0.3147110, -0.0902854, 0.0266519, -0.0611271, 0.0036804, 0.1580530, 0.0495644, -0.2001100, -0.1285720, -0.0125825, -0.0050515, 0.0005593, 0.0002059, -0.0000869, -0.0010948, -0.0028433, 0.1390820, 0.1378640, 0.1368050, 0.1427460, -0.2829230, -0.3412290, -0.4193620, -0.2941600, -0.1697150, -0.3723930, -0.1872180, -0.1696730, -0.2390840, -0.0509064, -0.0778084, -0.0036506, 0.1580000, 0.1043160, -0.0308885, -0.0929112, 0.0106104, -0.0247032, 0.0054019, 0.0004177, -0.0002430, 0.0003562, -0.0005988, 0.0009260, 0.1406170, 0.2896950, 0.1978670, 0.1061990, 0.0235411, -0.0898917, -0.2491810, -0.1347800, -0.3191410, -0.3287450, -0.2371600, -0.1219750, -0.0676829, -0.0352835, -0.0401429, 0.0063719, 0.0813171, 0.0333668, -0.2176720, -0.0934866, 0.0569034, -0.0408980, 0.0209995, 0.0012315, 0.0003614, 0.0005104, 0.0040417, 0.0096647, 0.1432340, 0.2453870, 0.1498210, 0.1583340, 0.2263560, -0.0640398, -0.0385070, -0.1729210, -0.2318350, -0.1397470, -0.3255070, -0.2921090, -0.1064310, 0.0948562, 0.0759362, -0.0134470, 0.2519160, 0.0091840, -0.2037610, -0.2015150, 0.0642170, -0.0234020, 0.0190314, 0.0057835, -0.0002004, 0.0006386, 0.0088430, 0.0525382, 0.0692433, 0.2401630, 0.2036420, 0.2097750, 0.2271810, 0.0090197, 0.2889710, -0.0348080, -0.0872451, -0.0992461, -0.2614590, -0.0274472, 0.1100150, 0.1806880, 0.0854857, -0.0186297, -0.1288730, -0.1561720, -0.0788465, -0.2096180, 0.0197370, 0.0628338, 0.0163877, 0.0146900, -0.0000704, 0.0002822, 0.0072169, 0.0982001, 0.0804236, 0.1784220, 0.0808836, 0.0726873, 0.1726680, 0.1789890, 0.4068810, 0.3051860, 0.0133914, -0.1707440, -0.1428970, 0.1191970, 0.1517050, 0.1177700, 0.1801700, 0.1166880, -0.0248936, -0.0259913, 0.1339540, -0.0351275, 0.0547384, 0.0677410, 0.0091956, 0.0030416, 0.0003171, -0.0004694, -0.0130718, 0.0583364, 0.0904228, 0.1469020, 0.0624813, 0.1503480, 0.1572850, -0.0104282, 0.2127490, 0.1192730, 0.3248350, 0.2220090, -0.0163725, 0.1217600, 0.1835000, 0.0233312, 0.1913170, 0.1368730, 0.1544590, -0.0390640, 0.0005818, 0.0225376, 0.0183991, 0.0360541, 0.0078093, 0.0012602, -0.0003145, -0.0012485, -0.0150858, 0.0654054, 0.0665722, 0.1239580, 0.0767589, -0.1077210, -0.0053320, 0.0507034, 0.0728776, 0.0779390, 0.0204226, -0.2118690, -0.1626220, -0.0479760, 0.2380400, 0.0563930, -0.0308087, 0.2076110, 0.1236530, 0.0568596, 0.1090240, 0.1543630, 0.1443590, 0.0378969, 0.0029602, 0.0006969, 0.0001401, -0.0000540, 0.0020182, 0.0188934, -0.0485785, -0.1066260, -0.0895276, -0.0275116, -0.0385695, -0.0590843, -0.0409029, -0.0396031, -0.0708542, -0.0435234, -0.0277954, 0.0707455, 0.1473840, -0.0129485, 0.0113855, 0.1758400, 0.2077500, 0.2228510, 0.3021800, 0.2455880, 0.1472850, 0.0254451, 0.0040501, -0.0007483, 0.0002755, 0.0002169, 0.0020780, -0.0216156, -0.1166020, -0.1168000, -0.0799220, -0.0365556, 0.1370460, 0.2976510, -0.1154210, -0.0173727, 0.0908094, 0.0148827, -0.0046308, 0.0352125, 0.0574678, -0.0065793, 0.1686000, 0.0281411, 0.1914500, 0.3631830, 0.3547160, 0.1496470, 0.0966839, 0.0102705, -0.0005999, 0.0005387, 0.0000975, -0.0002297, -0.0003617, -0.0067530, -0.1344970, -0.0905923, 0.0799211, 0.0106485, -0.0773186, -0.0646803, -0.0564052, 0.2151190, 0.1445770, -0.0868904, -0.0573881, -0.1274600, -0.1515030, 0.1525580, 0.2343620, -0.0137595, 0.0588639, 0.1777300, 0.1464320, 0.0689518, 0.0779366, 0.0137410, -0.0005211, -0.0000753, 0.0002275, -0.0001325, -0.0040152, -0.0058660, -0.0030172, -0.0131891, 0.1036820, 0.0915589, -0.0350359, -0.0566994, -0.2923160, -0.2187150, 0.0099168, -0.0515647, 0.0225287, -0.0507387, -0.0292343, 0.1643190, 0.1319620, -0.0426105, 0.0341211, 0.0882131, 0.1273560, 0.0452964, 0.0291230, 0.0111251, 0.0027703, 0.0000182, -0.0003117, -0.0006764, -0.0001513, 0.0018288, 0.0342891, 0.0728698, 0.0574413, -0.0018842, -0.1061150, -0.1180560, -0.0459243, 0.0642005, 0.0079470, -0.0805064, -0.0906607, -0.1744180, -0.1233070, -0.0143498, 0.0293696, 0.0258253, 0.0612719, 0.0523061, 0.0301489, 0.0003133, 0.0025752, 0.0028165, 0.0034401, -0.0001062, 0.0004196, 0.0000774, -0.0002161, -0.0001728, 0.0081637, 0.0503565, 0.0750133, 0.0286757, -0.0157914, -0.0509397, -0.0260569, -0.0473439, -0.0556514, -0.0832980, -0.0844420, -0.0914444, -0.0660521, -0.0414272, -0.0003561, 0.0009492, 0.0084314, 0.0148603, 0.0153494, 0.0012203, 0.0006943, 0.0000833, 0.0001511, -0.0001569, -0.0003772, -0.0004881, 0.0002536, 0.0000278, 0.0001803, -0.0008143, -0.0013117, 0.0009273, 0.0008789, -0.0035291, -0.0047016, -0.0053119, -0.0063116, -0.0035364, -0.0069562, -0.0088573, -0.0056592, -0.0001286, 0.0090698, 0.0005639, -0.0008751, 0.0001927, 0.0012868, -0.0009867, -0.0002552, -0.0000611, 0.0000878, -0.0008361, -0.0002587, 0.0001746, 0.0006481, -0.0000320, -0.0007150, -0.0002747, 0.0002555, 0.0001745, 0.0005303, -0.0000804, 0.0003975, -0.0003843, 0.0004174, -0.0000157, -0.0000765, 0.0000834, 0.0004285, 0.0002994, 0.0003843, 0.0000129, -0.0001972, -0.0002326, 0.0001824, 0.0008242, 0.0004683, 0.0000247, -0.0002380, 0.0002741, -0.0002435, 0.0002482, -0.0002733, 0.0005891, 0.0002853, 0.0006946, 0.0001132, 0.0002043, -0.0011092, -0.0011895, -0.0003888, 0.0005579, 0.0055768, 0.0057624, 0.0073438, 0.0199549, 0.0210336, 0.0099152, 0.0039974, 0.0043774, 0.0028602, 0.0052886, 0.0006740, -0.0001331, 0.0000862, 0.0004232, -0.0000030, -0.0004679, -0.0007525, -0.0003504, 0.0002465, -0.0000424, 0.0004444, -0.0003057, -0.0003240, 0.0019891, -0.0055015, -0.0232258, -0.0351598, -0.0190397, 0.0002478, -0.0017703, -0.0085884, -0.0267754, -0.0386917, 0.0197357, 0.0148432, 0.0391995, -0.0213753, -0.0171038, -0.0020313, -0.0029284, -0.0021974, -0.0002891, 0.0001233, -0.0005369, -0.0000081, -0.0001679, -0.0006055, -0.0002479, 0.0010899, 0.0021008, 0.0030285, -0.0117212, -0.0419867, -0.0503524, -0.0312044, -0.1011330, -0.0427528, -0.0668804, -0.0617702, 0.0111532, 0.0214485, 0.0086347, 0.0358447, 0.1795310, 0.1482100, 0.0421356, -0.0187262, -0.0250910, 0.0105858, -0.0010128, -0.0002122, 0.0002071, -0.0000957, -0.0001585, -0.0008102, -0.0001512, -0.0012626, -0.0046876, -0.0328541, -0.0499690, -0.0639136, -0.0817277, -0.0481895, -0.1111510, -0.0321568, -0.0204351, -0.0123563, 0.2533740, 0.1268790, 0.0159760, 0.0044251, 0.1222040, 0.0846725, 0.0762629, -0.0815391, -0.0229973, -0.0067159, 0.0154469, -0.0054720, -0.0003641, -0.0006883, -0.0001048, -0.0016104, -0.0062649, -0.0354207, 0.0179850, 0.0750067, 0.0625679, -0.0093240, -0.0194738, 0.0052780, -0.0778006, 0.0098282, 0.1279560, 0.1645100, 0.1790090, 0.2285180, 0.3492730, -0.0654064, -0.2910290, -0.0150815, 0.0738833, 0.0554411, 0.1273020, 0.0310634, -0.0666249, 0.0025767, -0.0001727, -0.0003507, -0.0000816, -0.0004990, -0.0458494, -0.0269906, 0.0862817, 0.1348890, 0.0352288, 0.0018804, -0.1680970, -0.0271150, 0.0741148, 0.0008800, 0.0906127, 0.1337920, -0.0081554, 0.2504280, 0.0715212, 0.0193170, -0.1932540, -0.2272060, -0.0260486, 0.0664388, 0.0291418, 0.1462910, 0.0739487, 0.0408274, 0.0030597, -0.0000547, -0.0007469, -0.0060810, -0.0518455, -0.0111431, 0.1150160, 0.0285120, -0.0286129, -0.1264900, 0.0395266, 0.0632243, 0.0231511, -0.0566849, 0.1022930, 0.2697380, 0.0683115, 0.4295320, 0.2720100, -0.0986501, -0.0867964, -0.0976981, -0.2172350, -0.0378465, 0.0562545, 0.0910191, 0.0964885, 0.0776640, 0.0001599, 0.0005195, 0.0022636, -0.0093953, -0.0160254, -0.0033596, 0.0352158, -0.1786110, -0.1868440, -0.0736730, 0.1686840, 0.0362285, -0.0487038, 0.2183960, 0.0166699, -0.0887319, 0.3959540, 0.2262130, 0.0205983, -0.2080710, -0.4019070, 0.0149047, -0.1130200, -0.0244812, 0.0674098, 0.2990900, 0.1895970, 0.0495423, -0.0027480, -0.0003620, 0.0015558, 0.0093289, -0.0182547, 0.0258218, -0.0712324, 0.0152798, 0.1111170, -0.0111364, -0.0494013, -0.0483949, -0.0009599, 0.1418150, -0.0186881, 0.5532970, 0.8211160, 0.1512240, -0.2881140, -0.1845810, -0.3788870, -0.2247120, -0.1296290, -0.0819578, 0.1790130, 0.2899370, 0.1784340, 0.0489426, 0.0299286, -0.0006350, 0.0009361, 0.0083442, -0.0204604, -0.1130470, -0.0945063, 0.1122270, -0.0509775, -0.2682610, -0.0918914, -0.0988056, -0.0504850, 0.1314350, 0.3339780, 0.7488780, 0.6120310, -0.0691230, -0.3999120, -0.4360930, -0.4027480, -0.2807990, -0.2163330, -0.2242370, -0.0396149, 0.2272640, 0.2892270, 0.0736477, 0.0072853, 0.0003151, 0.0006926, -0.0051681, 0.0097771, -0.1468390, -0.0172964, 0.1408750, -0.2646290, -0.2214250, -0.2076570, 0.0339760, 0.1940880, 0.2036980, 0.3499330, 0.4406230, -0.0847823, -0.6811930, -0.6908620, -0.4342870, -0.4032610, -0.4535740, -0.4141250, -0.3728650, -0.1253370, 0.0164411, 0.1194170, 0.0066170, 0.0013737, 0.0006502, -0.0007027, 0.0009598, 0.0567924, -0.1079120, -0.1062080, 0.1019670, -0.0574271, 0.0173319, 0.0604951, 0.1502090, 0.2264160, 0.4020120, 0.4102350, 0.1851850, -0.4810530, -0.6394770, -0.4802470, -0.2388800, -0.3982730, -0.3072730, -0.5108000, -0.3402290, -0.1489640, -0.0788200, 0.0213104, 0.0224818, -0.0016851, 0.0012056, -0.0014892, 0.0004271, 0.0463073, -0.0518246, -0.0670857, -0.0298271, 0.2037400, 0.0232724, 0.2269460, 0.3570100, 0.1759020, 0.2082280, -0.0279224, -0.1845210, -0.4577220, -0.2186160, -0.0958769, -0.2483690, -0.3979040, -0.3793170, -0.3479400, -0.4212560, -0.1375540, 0.0335348, -0.0014797, -0.0091795, -0.0077587, 0.0007658, -0.0010925, 0.0013582, 0.0118982, 0.0566331, 0.0122866, -0.0253047, 0.0172422, 0.0364255, 0.1908920, 0.1575360, 0.0352299, 0.0663503, -0.2286240, -0.3693630, -0.3338670, -0.2752030, -0.3326570, -0.2206130, -0.3285370, -0.2408310, -0.1645060, -0.1132340, -0.0115440, 0.1992560, -0.0064573, -0.0156673, -0.0010314, 0.0006118, 0.0001056, 0.0025116, -0.0030425, 0.0931030, 0.1188890, 0.0161423, 0.1050660, -0.0019846, 0.1869960, 0.0318862, 0.0056512, 0.1032060, -0.1124510, -0.3276760, -0.4297360, -0.3761720, -0.1535510, -0.1177850, -0.2494940, -0.2098620, -0.0481124, 0.0683082, 0.2717050, 0.2375760, -0.0330297, -0.0037631, -0.0016102, -0.0010583, -0.0000128, 0.0031463, -0.0011572, 0.0340262, 0.0153869, -0.0366232, -0.0764299, 0.1054450, 0.1401550, -0.0478824, -0.1284320, -0.0967892, -0.4176340, -0.3012060, -0.1795050, -0.1680250, -0.2213710, -0.1172750, 0.0686823, 0.1911500, 0.1276300, 0.1528730, 0.3299200, 0.1976660, -0.0582059, -0.0349747, -0.0004854, -0.0003291, -0.0002268, 0.0072013, 0.0440731, 0.0349688, 0.0568590, 0.0359108, 0.0263035, 0.1043590, 0.0875935, 0.0817035, 0.1639450, -0.2054030, -0.3443350, -0.1733930, -0.0919708, -0.0883710, 0.0305653, 0.1251720, 0.1886730, 0.0927039, 0.1126550, 0.3338860, 0.2971710, 0.1375810, -0.0171058, -0.0091200, -0.0039726, -0.0025421, 0.0001628, -0.0059057, 0.0368439, 0.1110000, 0.1466340, 0.0993838, 0.1479440, 0.0885706, 0.0836699, 0.1247540, 0.0399075, -0.1530670, -0.3075990, -0.1350360, -0.0020985, 0.1578460, 0.1023510, 0.1747230, 0.0848397, 0.3157670, 0.1793910, 0.2627050, 0.1954640, 0.0369550, 0.0027559, -0.0037975, 0.0044226, -0.0004784, 0.0010119, -0.0023652, 0.0037578, 0.0822302, 0.1289460, 0.1204940, -0.0171371, -0.1760750, -0.1581080, -0.0069986, 0.0202567, 0.1291490, -0.0179799, -0.0508358, -0.0028012, 0.1830190, 0.0141987, 0.2435770, 0.0925438, 0.3092330, 0.1817170, 0.0989350, 0.0145372, 0.0470134, 0.0338207, -0.0042355, 0.0028108, 0.0005765, 0.0012536, -0.0045593, -0.0613747, 0.0086269, 0.0828847, 0.0613850, -0.0852318, 0.0905872, 0.1273790, 0.1016560, 0.0301361, 0.1479810, 0.0837919, 0.0755858, -0.0563676, 0.0586855, 0.1531980, 0.2388640, 0.1955630, 0.1411650, 0.1213920, -0.0138424, 0.0207818, 0.0234921, 0.0245456, -0.0011928, 0.0007086, -0.0001567, -0.0010327, -0.0226007, -0.0825733, -0.0591471, -0.0016505, -0.0410770, -0.1364060, -0.0857768, -0.1584180, -0.0769056, -0.0520954, 0.1751850, 0.0368436, 0.0033223, 0.1301450, 0.0300255, -0.0418817, 0.0883899, 0.0586992, 0.0970506, 0.0702717, -0.0203448, 0.0093890, 0.0210116, 0.0732231, 0.0030843, 0.0002907, 0.0003453, -0.0000394, -0.0091681, 0.0127650, -0.0098256, 0.0052565, -0.0701238, -0.0414344, -0.0638839, -0.0001040, -0.0395935, 0.0553929, 0.1022450, 0.1388510, 0.0423214, 0.1869270, 0.0125729, 0.0714369, 0.1314390, 0.0764887, -0.0464743, -0.0340287, 0.0088723, -0.0344228, 0.0112902, 0.0340725, 0.0143632, 0.0000212, -0.0003960, 0.0000335, -0.0012004, 0.0268143, 0.0997296, 0.1068610, 0.0258992, -0.1844310, -0.1001750, 0.1055090, 0.1040250, -0.1397130, -0.0653816, -0.0036200, 0.1501880, -0.0165623, -0.0157449, 0.1479480, 0.0871873, 0.1422950, -0.0094228, -0.0842706, -0.0792720, -0.0183119, 0.0038813, 0.0376272, 0.0120458, -0.0000700, -0.0002397, -0.0006005, -0.0001993, -0.0002597, -0.0081898, 0.0476529, 0.0244242, 0.0897341, 0.0111093, 0.1882040, 0.1173010, 0.0115902, 0.0520154, -0.0364249, 0.0250169, 0.0575586, -0.1013380, 0.1927980, 0.1028830, 0.0723711, 0.0040776, -0.0275897, -0.0398080, -0.0516613, -0.0124905, -0.0066755, 0.0005023, 0.0000682, 0.0001384, -0.0001691, -0.0002460, 0.0008499, -0.0031065, -0.0274522, -0.0773880, -0.0207319, -0.0654206, 0.0376162, -0.0608794, 0.0502546, 0.1638970, 0.0698406, -0.1347650, -0.1574340, -0.1456830, -0.0202549, -0.0162161, 0.0099243, 0.0082133, -0.0441146, 0.0386748, 0.0140405, 0.0068779, 0.0004355, 0.0000326, -0.0002612, -0.0000028, 0.0006267, -0.0000732, -0.0003186, -0.0010277, -0.0225015, -0.0560590, -0.0648570, -0.0617670, -0.0460139, 0.0007752, -0.0087953, 0.0275937, -0.0393306, -0.1072630, -0.0431816, -0.0275952, -0.0828701, -0.0409883, 0.0357058, -0.0420004, -0.1200110, -0.0296154, -0.0027487, -0.0013417, -0.0000452, 0.0005877, 0.0002829, -0.0001448, -0.0000496, -0.0000772, -0.0004530, 0.0000564, -0.0001566, -0.0006553, -0.0089258, -0.0094504, -0.0012844, 0.0011942, -0.0044040, -0.0125103, -0.0184731, -0.0321372, -0.0537890, -0.0217715, -0.0161974, -0.0347120, -0.0087354, -0.0067729, -0.0425289, -0.0325502, -0.0014110, -0.0002970, 0.0005677, -0.0003756, -0.0007236, 0.0002801, 0.0002389, 0.0003999, -0.0000245, -0.0002774, -0.0001879, -0.0001566, 0.0000429, -0.0000287, 0.0002847, 0.0002369, -0.0001759, -0.0004662, 0.0002570, 0.0000999, 0.0007131, -0.0000115, -0.0001577, 0.0005232, -0.0000683, -0.0000068, -0.0000419, -0.0004304, 0.0001840, -0.0001278, 0.0001436, -0.0002830, 0.0007245, 0.0001889, -0.0000100, 0.0001419, -0.0006031, -0.0001853, 0.0001037, 0.0002769, -0.0004021, 0.0006647, 0.0014942, 0.0042021, 0.0027012, 0.0003503, 0.0008272, 0.0011765, 0.0136629, 0.0029592, -0.0001154, 0.0002950, 0.0012119, 0.0047489, 0.0019625, 0.0001575, 0.0007824, 0.0002195, 0.0000935, -0.0000641, 0.0000122, 0.0002737, -0.0007158, -0.0002899, 0.0004179, -0.0006065, -0.0003556, -0.0014035, 0.0003214, -0.0004576, 0.0000243, 0.0111622, 0.0060258, -0.0062869, 0.0179304, 0.0576656, 0.1181090, 0.0924536, 0.0366394, 0.0217068, 0.0159953, 0.0041021, -0.0005517, -0.0000080, -0.0000559, -0.0001629, 0.0001569, 0.0002195, -0.0004043, -0.0000556, 0.0001065, 0.0002143, -0.0001797, 0.0007231, 0.0282681, 0.0242430, 0.0320123, 0.0520214, 0.0074905, 0.0624408, 0.1151440, 0.1394600, 0.2446320, 0.3135380, 0.1822450, 0.1280990, 0.1870390, 0.1784240, 0.1031770, 0.1363960, 0.0581387, -0.0018080, -0.0109534, -0.0009986, 0.0005159, 0.0002448, 0.0001488, 0.0000910, 0.0000088, -0.0019537, 0.0008002, 0.0053868, 0.0226831, -0.0100613, 0.0144678, 0.0454928, 0.0853818, 0.1900570, 0.3480730, 0.3626690, 0.2348640, 0.1620940, 0.1899840, -0.0306146, -0.2242020, -0.0763052, -0.0445284, -0.0509790, 0.0216416, 0.0231297, 0.0292506, 0.0023595, -0.0004371, -0.0035911, -0.0009730, 0.0003784, 0.0000489, -0.0000983, 0.0142760, 0.0192135, 0.0522465, 0.0444215, -0.0098425, -0.0298511, 0.0901989, 0.2211860, 0.1466830, 0.0165682, 0.0220348, 0.0475385, 0.0742537, -0.0969036, -0.0065055, 0.0345777, 0.0363538, -0.0005766, -0.0749331, 0.0091792, 0.0215467, -0.0306701, -0.0124163, -0.0041694, -0.0015915, 0.0003078, 0.0004276, 0.0067798, -0.0436115, -0.0517953, -0.1080000, -0.0635494, 0.0144669, -0.0511079, 0.0357250, 0.0602577, 0.0482169, -0.0608304, -0.0156686, 0.1404020, 0.1836140, 0.2174850, 0.0341271, 0.1053450, 0.1896220, 0.1236570, -0.0386304, 0.0962878, 0.0419897, -0.0351545, -0.0218656, 0.0218132, -0.0018379, 0.0002771, -0.0028205, -0.0069702, -0.0487734, -0.1017230, -0.1220450, 0.0229833, -0.1657720, -0.0859261, 0.1766410, 0.3160120, 0.3440200, 0.1463020, 0.0614506, 0.1222740, 0.0407970, 0.0525580, 0.1731980, -0.0746411, 0.0934179, 0.1005630, -0.1364170, 0.0518141, -0.0217160, 0.0206613, 0.0275086, 0.0233224, 0.0001459, 0.0030362, -0.0129674, -0.0269569, -0.0158916, -0.1975320, -0.0503149, -0.0041884, -0.2863320, -0.1021320, 0.1656560, -0.0261896, 0.0670890, -0.0052077, 0.0451364, 0.2279320, 0.1428580, -0.0440824, 0.0211099, 0.1365890, 0.0402627, -0.1487490, -0.0125310, -0.0368251, -0.2132100, -0.0528429, 0.0475223, -0.0022897, 0.0009809, -0.0002179, -0.0155109, -0.0230223, -0.0430363, -0.1508780, -0.1215720, 0.0480891, -0.1293020, -0.1992690, 0.0656448, -0.0672274, 0.0683811, 0.0262810, -0.0673850, -0.1858980, -0.1099450, 0.0517338, 0.0441837, 0.1327910, 0.0805458, -0.0023643, -0.0377358, 0.0033369, -0.2575700, -0.0443654, -0.0272144, -0.0528958, -0.0059388, 0.0002671, -0.0145693, -0.0349260, -0.0457083, -0.1666200, -0.1221910, -0.0194230, -0.0068186, 0.0410390, 0.0782512, -0.1721530, -0.0241591, 0.0426622, -0.2480890, 0.0779159, -0.0092481, 0.0932035, 0.0933988, 0.0128376, 0.0327752, -0.0514601, -0.1752630, -0.0343052, -0.0949660, -0.0965098, 0.0257076, -0.0300853, -0.0034702, -0.0001797, -0.0110976, -0.0854488, -0.1341980, -0.2481960, -0.2614280, -0.2052560, -0.2705900, -0.0611990, -0.2724430, -0.1706110, -0.1333100, -0.0588962, 0.1188120, 0.2276320, -0.0160405, -0.1007990, 0.1542850, 0.1257610, -0.1846850, -0.1298860, -0.0071449, 0.1455320, -0.0137841, -0.0330909, 0.0192708, -0.0283488, 0.0001045, -0.0003550, -0.0052919, -0.0717785, -0.2114600, -0.2045260, -0.3405200, -0.1786310, -0.4253450, -0.3521220, -0.3347990, -0.0196060, 0.2194250, 0.2325770, 0.3693290, 0.2065130, 0.1604280, 0.1217200, 0.1145720, 0.0782240, -0.1677220, -0.1115720, -0.0118817, 0.1478640, 0.1526960, -0.0607611, -0.0214455, 0.0010462, -0.0012636, 0.0001006, -0.0029469, -0.0570988, -0.1652610, -0.1496500, -0.2126220, -0.2810670, -0.0527090, -0.0509214, -0.2104870, 0.0629435, 0.2724750, 0.6655810, 0.2977940, 0.0317322, 0.2046410, 0.2998310, 0.1067240, -0.0517592, 0.2841260, 0.0221685, 0.1293210, 0.0127886, 0.2382930, 0.1381650, 0.0089277, -0.0016301, -0.0009651, -0.0004155, -0.0013186, -0.0332156, -0.0618432, -0.0609062, -0.0972372, -0.0288386, -0.0084770, -0.0476495, 0.2624420, 0.4386990, 0.8190360, 0.5641870, 0.0294079, -0.2326160, 0.1235190, 0.3611170, 0.2262860, 0.1548350, 0.1360620, 0.3326090, 0.0977511, 0.1531500, 0.2414780, 0.1701020, 0.0277205, -0.0029329, -0.0000284, 0.0004865, 0.0029950, -0.0032807, -0.0277997, 0.0939376, 0.1582750, 0.1766970, 0.0471980, 0.3750710, 0.5056110, 0.7608620, 0.5279880, 0.1178220, -0.2540620, -0.1969960, 0.1063300, 0.3318890, 0.3282210, 0.3453460, 0.2849970, 0.2433110, 0.2830210, 0.1612170, 0.1364630, 0.0450439, 0.0154647, -0.0064892, -0.0066415, 0.0003898, 0.0013484, 0.0024170, -0.0270397, 0.1629060, 0.3864260, 0.3214300, 0.4378460, 0.6549810, 0.7692930, 0.6037570, 0.1829690, -0.1707280, -0.3602500, -0.0058983, -0.0226519, -0.2991550, 0.0269918, 0.1279340, 0.0470282, 0.2502260, 0.1572330, 0.2332690, 0.0725069, 0.0246352, -0.0380436, -0.0239080, -0.0129137, 0.0002055, 0.0006964, -0.0005722, 0.0048549, 0.1618020, 0.3405300, 0.5088260, 0.8238170, 0.9051550, 0.7926690, 0.2607440, -0.1724900, -0.4467350, -0.2878370, -0.1854990, 0.0142654, -0.1712420, -0.2773960, -0.0890615, -0.0318082, -0.0155739, -0.0498147, 0.1558440, 0.1072870, 0.0306810, -0.0443087, 0.0026366, -0.0019475, -0.0002893, 0.0001410, -0.0033740, 0.0172207, 0.1158850, 0.2831830, 0.4732930, 0.6339380, 0.6033350, 0.2225800, -0.0901998, -0.2179170, -0.3956850, -0.3252840, -0.1715190, -0.2603230, -0.0021407, 0.0097198, -0.1522820, -0.0022263, 0.0060270, 0.0640781, 0.1100070, 0.1041110, -0.0101735, -0.0340286, -0.0059340, -0.0013647, -0.0001604, -0.0035676, -0.0083348, 0.0550610, 0.0798368, 0.2752450, 0.3941450, 0.4164600, 0.1968520, -0.1560650, -0.2401600, -0.4441770, -0.1947920, -0.4466490, -0.3350530, -0.1246320, 0.0331608, -0.0777392, -0.0506659, 0.0659314, -0.0273174, 0.1337360, 0.1263620, 0.0220522, -0.0195867, -0.0352314, -0.0072516, -0.0000854, 0.0002527, -0.0002052, -0.0145561, -0.0210547, 0.1290850, 0.2638820, 0.2753240, 0.1965060, 0.0331011, -0.0454606, -0.1735030, -0.3526500, -0.3506750, -0.0384169, -0.1069150, -0.3079420, 0.0440772, -0.0544711, -0.0623159, 0.0317376, -0.0822028, -0.0800045, 0.0208689, -0.0197318, -0.0185956, -0.0339520, -0.0044389, 0.0004303, -0.0003318, 0.0000352, -0.0187588, -0.0329108, 0.1455080, 0.1637180, 0.0704819, 0.1470340, 0.0962120, 0.1242090, -0.1502650, -0.1383810, -0.1379110, -0.0926272, -0.2083870, -0.3324890, -0.1106940, -0.2504390, -0.1154610, -0.2376970, -0.1536680, -0.1382130, -0.0282946, -0.0356829, -0.0050114, -0.0293286, -0.0034205, -0.0003726, -0.0006819, 0.0001569, -0.0060951, 0.0120291, 0.0501300, -0.0273715, -0.0854135, -0.1459760, -0.1445320, -0.1153140, -0.0262309, -0.2301710, -0.1330930, -0.1169580, -0.1996380, -0.1398690, -0.0030776, -0.2621050, -0.1900920, -0.1916570, -0.0536675, -0.0655983, 0.0726907, -0.0211169, -0.0056225, -0.0157196, -0.0010825, -0.0002261, 0.0006297, -0.0006872, 0.0083768, 0.0573151, -0.0029269, 0.0424520, -0.0715130, -0.1307460, -0.1118570, -0.1351210, 0.0359885, -0.0385180, -0.1850700, -0.2590930, -0.0974517, -0.1847360, -0.3484020, -0.2491570, -0.1374210, -0.1665780, -0.0504818, 0.0334396, 0.0039366, -0.0396886, -0.0100811, -0.0067774, -0.0008111, -0.0000581, 0.0002102, 0.0005219, 0.0132525, 0.0344627, 0.0294862, 0.1084610, 0.1420160, 0.3240620, 0.1915770, 0.1347440, 0.0592767, -0.0439766, -0.1217000, -0.1791250, -0.1628430, -0.0312518, -0.0144072, -0.1053010, -0.1898320, -0.2573440, -0.0474896, -0.0079453, -0.0242568, 0.0146859, -0.0080687, -0.0033524, -0.0004640, -0.0000155, -0.0000563, -0.0001441, 0.0028656, -0.0058796, 0.0056901, 0.0949191, 0.0007419, 0.0664681, 0.1210740, 0.1602540, 0.1947410, 0.1479530, -0.0090073, 0.0741906, -0.0251016, -0.1891740, -0.0063987, -0.1369150, -0.0785071, -0.0269018, 0.0109657, 0.0143215, -0.0073961, 0.0085344, 0.0023289, 0.0009721, 0.0002622, -0.0002885, 0.0005520, -0.0005560, 0.0001268, 0.0000831, 0.0214011, 0.0654145, 0.0770458, 0.0494813, -0.0021396, 0.0148340, 0.0500091, 0.0767832, 0.1132600, 0.0290508, 0.1279150, 0.1348160, 0.1193420, 0.0758383, 0.0618851, -0.0709092, -0.0281355, 0.0343764, 0.0038560, 0.0005806, 0.0003313, -0.0004386, 0.0005839, 0.0000802, -0.0003558, -0.0002594, -0.0001263, 0.0002220, -0.0001142, -0.0007534, -0.0017103, -0.0035062, -0.0056984, -0.0159673, -0.0387859, -0.0015057, -0.0033972, -0.0561481, -0.0127286, 0.0692485, 0.0034327, 0.0038574, 0.0811692, -0.0045304, 0.0005554, 0.0097313, 0.0102914, -0.0005889, 0.0005645, -0.0000031, -0.0001730, -0.0001614, -0.0005667, 0.0006230, 0.0006882, -0.0005658, -0.0002933, 0.0004173, 0.0002995, 0.0000346, -0.0001986, 0.0000808, -0.0003399, -0.0000684, 0.0000797, -0.0000814, 0.0002895, -0.0010995, 0.0001200, 0.0000084, -0.0005843, -0.0002701, -0.0000881, 0.0001134, -0.0001260, 0.0003366, 0.0006167, 0.0006678, -0.0000554, 0.0004189, 0.0000893, -0.0000224, -0.0004049, 0.0008025, 0.0001111, 0.0004475, -0.0000216, -0.0002089, -0.0004898, -0.0012239, -0.0058355, -0.0050738, -0.0004691, 0.0000818, -0.0010610, -0.0024087, -0.0029529, -0.0010587, -0.0007563, -0.0002573, -0.0000465, 0.0001707, 0.0003913, 0.0001207, -0.0002230, -0.0002591, 0.0002238, 0.0002661, -0.0000714, -0.0003441, -0.0004538, 0.0000895, 0.0002042, -0.0004505, -0.0085030, -0.0083119, -0.0127296, -0.0227340, -0.0268591, -0.0229570, -0.0292380, -0.0289563, -0.0393646, -0.0399352, -0.0252294, -0.0093348, -0.0249446, -0.0122459, -0.0077826, -0.0003035, 0.0015907, -0.0013293, -0.0001661, -0.0000918, -0.0000506, -0.0001915, 0.0004414, 0.0002290, 0.0001993, -0.0020942, -0.0122819, -0.0052984, -0.0164936, -0.0259897, -0.0420660, -0.0578622, -0.0600867, -0.0237356, 0.0276175, 0.0737825, 0.0703193, 0.0194550, 0.1067560, 0.0946741, -0.0190245, -0.0187709, 0.0011252, -0.0149643, -0.0008711, 0.0008134, -0.0012121, 0.0000544, -0.0003491, 0.0001820, 0.0003851, -0.0005758, 0.0003301, 0.0009222, -0.0037041, -0.0202733, -0.0282360, -0.0480622, -0.0567391, -0.0372964, -0.0463741, 0.0007000, 0.0133555, 0.0411253, 0.0422093, 0.0967127, 0.2033740, 0.2005330, 0.1527810, 0.1406810, 0.0457139, -0.0376777, 0.0161218, 0.0067341, -0.0281181, -0.0087725, -0.0041570, -0.0000511, 0.0004874, -0.0003158, 0.0003627, -0.0082304, 0.0005253, 0.0060748, 0.0016142, 0.0173191, 0.1555300, 0.1422700, 0.0140628, -0.2129900, -0.1148760, 0.0338063, -0.0431997, -0.2205090, -0.2019580, -0.0822662, 0.0171313, 0.0661130, 0.0574794, 0.0254291, 0.0210425, 0.0033605, -0.0389003, -0.0216970, -0.0095234, -0.0056531, 0.0003091, -0.0002007, 0.0052993, 0.0236999, 0.0607256, 0.0591163, -0.0222433, 0.0018385, 0.0933253, -0.1970270, -0.2413400, -0.0686592, 0.1731860, 0.2537860, -0.1374950, -0.3235470, -0.2379800, 0.0357461, 0.0726241, 0.0471046, -0.0276755, 0.1295310, 0.1013860, 0.0457077, -0.0317773, -0.0524889, -0.0341115, -0.0185260, -0.0003744, 0.0035907, 0.0136092, 0.0616321, 0.0326874, -0.0580055, -0.0009059, 0.1166010, -0.0077896, 0.1283830, 0.1754620, 0.0458934, 0.0640928, 0.1172480, -0.0837915, -0.3307850, -0.2689110, 0.0126440, 0.3099480, -0.0087194, -0.1758120, -0.1286500, -0.0094900, -0.0254977, -0.0675336, -0.0614813, -0.0352599, -0.0028377, 0.0108713, 0.0107563, 0.0452657, 0.0563960, -0.0169068, 0.0028538, -0.0251749, 0.0664252, 0.1513150, 0.0827030, 0.0955504, -0.0524579, 0.2424460, -0.0053148, 0.0048174, 0.0899591, -0.2616820, 0.0351130, 0.2346510, -0.1781660, 0.0113377, 0.0192679, 0.0778704, 0.1069870, -0.0317074, -0.0779012, -0.0367743, -0.0042676, 0.0006894, 0.0100550, 0.0020346, 0.0600258, 0.1645220, 0.0841214, 0.1983780, 0.2367180, 0.1440860, 0.0956184, 0.0903805, 0.0823487, 0.1788320, 0.4016010, 0.1775290, 0.0669578, -0.0830930, 0.2176380, 0.2385970, 0.0837045, 0.1336660, 0.2194100, 0.1765210, 0.2226820, 0.0546699, -0.0294381, -0.0633567, -0.0015198, 0.0004585, 0.0097845, 0.0376001, 0.0406640, 0.1041010, 0.0275967, -0.0377814, 0.0907499, 0.0375024, 0.0458511, 0.1842570, 0.3053370, 0.2806010, 0.2839670, -0.0560089, -0.3424430, -0.1535470, 0.2140300, 0.1733800, 0.3407890, 0.3573910, 0.2412330, 0.1904150, 0.1622270, 0.0524749, -0.0290833, -0.0424751, -0.0004584, -0.0000864, 0.0118789, 0.0362701, 0.0581338, -0.1345060, -0.0520511, 0.0627840, -0.0726471, -0.3336580, 0.1200510, 0.1084520, 0.3169670, 0.1499030, -0.2845610, -0.6013500, -0.5419910, -0.0435585, 0.2264010, 0.2103380, 0.1447120, 0.2035400, -0.0320261, -0.0740803, 0.0617151, 0.1009990, -0.0389069, -0.0050336, 0.0000931, 0.0002655, 0.0062526, 0.0245231, 0.0158146, -0.1761110, -0.0520149, -0.0252370, -0.0013482, -0.0028943, 0.0979313, 0.0997726, 0.2489680, 0.0663547, -0.5304400, -0.7983470, -0.4640510, 0.2212650, 0.1905770, 0.1402360, -0.1598180, 0.0278611, -0.0439055, 0.0945336, 0.0078006, 0.1260820, -0.0388457, -0.0137009, -0.0001178, -0.0003199, 0.0037127, 0.0366990, -0.0061127, -0.1349450, -0.1113290, 0.0308516, -0.0572095, 0.1533250, 0.0798402, 0.0936833, 0.2398340, -0.1447090, -0.7136880, -0.9452390, -0.6264670, -0.0077018, 0.0501075, -0.0528185, -0.2905370, -0.0625703, -0.0381845, 0.0037373, 0.0181560, 0.0906043, 0.0359188, -0.0076028, -0.0003017, 0.0001754, 0.0034366, 0.0325196, -0.0123479, -0.1572200, 0.2272830, 0.0988312, 0.1651540, 0.0818708, 0.0845658, 0.4192810, 0.1634690, -0.3924990, -0.9101120, -0.6665900, -0.3389910, -0.1595250, 0.0318111, -0.0844660, -0.1062650, -0.2524480, -0.1443570, -0.0307993, 0.2514440, 0.1275820, 0.0206761, -0.0015685, -0.0003266, -0.0000443, -0.0003936, 0.0145401, 0.0329486, -0.1342470, 0.2415750, 0.0740032, 0.4111360, 0.0175262, 0.0402233, 0.2803550, -0.2181000, -0.7375220, -0.7100590, -0.4264360, -0.3178340, -0.2250760, 0.0239102, -0.1510660, -0.1139820, -0.1699720, -0.0852494, 0.1778160, 0.2877080, 0.0979567, -0.0425954, -0.0143958, -0.0013930, 0.0001132, -0.0004124, 0.0017331, 0.0239677, 0.0584451, 0.0688535, -0.0148080, 0.1788740, 0.0523009, -0.0567062, 0.0599134, -0.4895350, -0.6935880, -0.4936680, -0.0244292, 0.1115140, -0.1612690, -0.0697063, -0.2112130, -0.0510502, -0.0020187, 0.2160210, 0.0951772, 0.1857220, 0.0679346, -0.1024920, -0.0289139, -0.0032956, 0.0000953, -0.0005167, 0.0069372, -0.0188143, 0.0851114, 0.1585910, -0.0117272, -0.0529824, -0.1135750, -0.1358070, -0.1009270, -0.4532320, -0.5300360, -0.2983080, 0.1051420, -0.1544870, -0.1977340, -0.1821660, 0.0327547, -0.1261320, 0.0349484, 0.1304750, 0.1464500, 0.1167940, 0.0241719, -0.0347537, -0.0091664, -0.0002364, 0.0030072, 0.0001906, 0.0067373, -0.0301676, -0.0327989, 0.0237404, 0.0055706, 0.0786919, -0.0361582, -0.1450630, -0.1622870, -0.3315530, -0.3209850, -0.1508770, 0.1064830, -0.0767744, 0.0504183, -0.0546063, 0.1947290, -0.1371810, 0.1051930, 0.2252290, 0.1013430, -0.0190214, -0.0572942, -0.0081157, -0.0022195, -0.0011580, -0.0001824, 0.0166257, 0.0025660, -0.0122469, 0.0270424, -0.0311941, 0.0849588, 0.0483363, -0.0592016, -0.2253770, -0.3300510, -0.3037720, -0.2982690, -0.1430030, 0.0547605, -0.0978472, -0.1242880, 0.2411210, 0.0289276, 0.0143114, 0.1601570, 0.0870574, -0.0453559, -0.1494030, -0.1005900, -0.0106906, -0.0071600, 0.0002951, -0.0002271, 0.0003362, 0.0044723, -0.0052501, -0.0187963, -0.0702138, -0.0682386, -0.0282859, -0.0688531, -0.1399540, 0.0643363, 0.0496339, 0.1401490, -0.1022950, 0.0978890, -0.0087350, -0.0640016, -0.0814111, -0.0715062, 0.0960835, -0.0925998, -0.0575806, -0.1395920, -0.1998540, -0.1283040, -0.0476248, -0.0020112, -0.0002621, 0.0003920, -0.0000353, 0.0168382, 0.0161128, -0.0348428, 0.0032839, -0.1431300, -0.2660470, -0.0947222, 0.0636938, 0.2893770, 0.3507080, 0.1261320, -0.0393091, -0.0015837, -0.0553281, 0.1067960, -0.1042050, -0.0332803, -0.0880625, -0.0972718, -0.0104190, -0.0930822, -0.1128030, -0.0261392, -0.0004665, 0.0031397, 0.0001013, -0.0005126, 0.0001187, 0.0171679, 0.0059600, -0.0462865, 0.0109883, 0.0373591, -0.0666979, 0.0571774, 0.2048910, 0.0557344, 0.2116950, -0.0066588, 0.1831670, -0.1866120, 0.1681910, 0.0177272, -0.0754749, 0.0844497, 0.0052784, -0.1640420, -0.0611787, -0.1097130, -0.1140620, -0.0468511, 0.0023344, 0.0022438, -0.0000791, -0.0005351, -0.0000986, -0.0137495, -0.0305069, -0.0482508, -0.0342508, 0.1024460, 0.1162410, -0.0531819, 0.0318271, -0.0598462, 0.0182881, -0.0043188, -0.0678652, -0.0559047, 0.0676302, 0.0326128, 0.1349740, 0.0091680, -0.0741844, -0.1891350, -0.0648773, -0.1534470, -0.0896172, -0.0314735, 0.0027058, 0.0004805, 0.0005267, 0.0003781, 0.0009438, -0.0173488, -0.0171945, 0.0035963, 0.0525147, 0.0988822, 0.1454090, 0.1291230, 0.0549478, 0.0583568, -0.1556560, -0.1714990, -0.0614726, -0.1414170, -0.0482823, -0.1405860, 0.0140555, -0.0794118, -0.0904048, -0.2207910, -0.0309892, -0.1055310, -0.0639501, -0.0091582, -0.0026717, 0.0001311, -0.0003772, 0.0000916, -0.0002905, -0.0047178, -0.0007447, 0.0036638, -0.0949134, -0.0732099, 0.0051217, 0.2089550, 0.1101080, -0.0626947, 0.0577999, 0.2206310, 0.1518630, 0.1057350, 0.0382641, 0.1057540, 0.0091614, -0.0449963, -0.0893440, -0.1198450, 0.0423149, -0.0282626, -0.0341732, -0.0017705, 0.0001057, -0.0004540, 0.0001497, 0.0000484, 0.0002978, -0.0000365, 0.0001980, -0.0099393, -0.1704850, -0.2000450, -0.0924874, -0.0446552, -0.0177084, -0.0835429, -0.1114380, -0.0461170, 0.1015120, 0.0370076, 0.1083620, 0.1025370, 0.0701047, 0.1382280, 0.1537790, 0.0068234, 0.0031471, 0.0308601, -0.0050071, -0.0003528, -0.0001996, -0.0000242, -0.0000947, 0.0000709, -0.0002584, -0.0002205, 0.0000412, 0.0005046, 0.0015745, 0.0028505, 0.0047459, 0.0070964, 0.0171701, 0.0344825, -0.0007377, 0.0107496, 0.0793209, 0.0512707, -0.0834081, 0.0010751, 0.0512893, 0.0323947, -0.0060317, 0.0104056, 0.0483730, 0.0404660, 0.0047554, 0.0001733, -0.0000807, 0.0001192, -0.0000306, -0.0002575, 0.0006506, -0.0000165, -0.0002341, -0.0000496, 0.0004781, -0.0000058, -0.0002339, 0.0002224, 0.0001027, 0.0000858, 0.0001458, -0.0001354, 0.0001983, -0.0004779, -0.0006395, -0.0000333, -0.0002778, 0.0001217, -0.0005429, -0.0007007, -0.0001490, 0.0004087, 0.0006021, 0.0000443, -0.0003497, -0.0001424, -0.0001452, 0.0001683, -0.0000051, 0.0001802, 0.0000584, 0.0002804, -0.0002636, 0.0006907, 0.0001726, 0.0004157, -0.0002268, 0.0000755, -0.0039620, -0.0007062, 0.0018037, 0.0038067, 0.0097205, -0.0073454, -0.0025766, 0.0015019, 0.0025829, 0.0027125, 0.0001372, 0.0002034, 0.0012401, 0.0001251, 0.0005706, 0.0000065, -0.0001030, -0.0002225, -0.0001728, 0.0002882, 0.0000025, -0.0005847, -0.0007164, -0.0024757, -0.0019893, -0.0154745, -0.0499606, -0.0481969, -0.0368186, -0.0180680, 0.0496697, 0.0294116, 0.0655088, 0.0911638, 0.0157516, -0.0034726, 0.0123863, 0.0045184, 0.0078256, 0.0098626, 0.0034975, -0.0083348, -0.0060748, 0.0004500, -0.0004047, -0.0000984, 0.0000637, -0.0011850, 0.0003758, -0.0029514, 0.0253462, 0.0218812, 0.0214773, -0.0192673, -0.1194950, -0.1307230, -0.1185080, -0.0457739, -0.0353985, -0.0230544, 0.0179207, -0.0304619, -0.0736281, -0.0275707, -0.0349636, -0.0272726, 0.0134181, 0.0542110, 0.0477666, 0.0187777, -0.0253956, -0.0050771, 0.0004406, 0.0003131, -0.0007197, -0.0026566, -0.0003336, 0.0066799, 0.0293641, -0.0066855, -0.0411485, -0.0139287, -0.1875720, -0.1587890, -0.2051590, -0.1875660, -0.0141997, 0.0569409, 0.0077873, 0.0123806, -0.1523440, -0.1270550, 0.0186801, 0.0563475, 0.0858892, 0.1079840, 0.0232713, -0.0820396, -0.0569638, -0.0142396, 0.0015294, 0.0000747, -0.0001207, -0.0001791, 0.0053418, 0.0219685, 0.0253315, -0.0267579, -0.0869293, -0.2742910, -0.3698510, -0.3463050, -0.3073380, -0.2863110, -0.2729460, -0.3450370, -0.1315810, -0.2175960, -0.1276400, -0.1443350, -0.0686121, -0.0755733, 0.0140253, 0.0052205, 0.0638188, -0.0151211, -0.0764432, -0.0071363, 0.0040091, 0.0002978, 0.0005757, 0.0010972, 0.0194255, 0.0438214, 0.0159256, -0.0226074, -0.1622730, -0.3534620, -0.2963800, -0.5043070, -0.3509940, -0.3122440, -0.1829280, -0.2370870, -0.1984120, -0.0443908, -0.1370920, -0.0610280, -0.1996170, -0.0244345, -0.1262830, -0.0797998, 0.0063664, -0.0112178, -0.0498274, -0.0122936, 0.0079221, -0.0000904, 0.0000502, -0.0134944, 0.0214930, 0.0649294, 0.0525453, 0.0253849, -0.0482600, -0.2254540, -0.2713710, -0.4301070, -0.3835270, -0.3292570, -0.3206330, -0.0520170, -0.1928330, -0.2418880, -0.2750030, -0.2934870, -0.2787060, -0.0960583, -0.1707890, -0.1608460, -0.0620376, -0.0287308, -0.0354655, -0.0108452, 0.0009061, -0.0003587, -0.0008456, -0.0030898, 0.0522707, 0.1128000, 0.0942720, 0.0970453, 0.0196227, -0.0585748, -0.2191370, -0.2990060, -0.4931810, -0.6417410, -0.4664040, -0.4018500, -0.3620670, -0.3600650, -0.2206090, -0.2632550, -0.1603070, -0.2588500, -0.0539371, -0.2483680, -0.2097650, -0.0729848, -0.0028883, 0.0004186, -0.0003737, -0.0003379, -0.0002345, 0.0080519, 0.0623047, 0.1378290, 0.1607930, 0.2951320, 0.3864590, 0.1823160, 0.0701550, 0.0022722, 0.0895867, -0.1029260, -0.2093300, -0.1612520, -0.1594350, -0.1178230, -0.2742310, -0.0791302, -0.0526830, -0.2303540, -0.1499850, -0.1667800, -0.1603470, -0.0426125, -0.0264369, -0.0041699, -0.0020626, 0.0000519, 0.0004395, 0.0070205, 0.0659730, 0.1497730, 0.2100960, 0.3356690, 0.4233120, 0.3808360, 0.4716420, 0.4489850, 0.4227260, 0.4661500, 0.2972020, 0.2579900, 0.1127820, 0.0015535, -0.0321578, 0.0650542, 0.0850094, -0.1181510, -0.0868842, -0.1473040, -0.0350349, -0.0158135, -0.0544760, -0.0194352, -0.0005595, 0.0006765, -0.0013746, 0.0117913, 0.0531959, 0.1480960, 0.2386570, 0.2355140, 0.2455400, 0.4078880, 0.4903960, 0.3618320, 0.1617860, 0.2159180, 0.4014690, 0.2457620, 0.3551910, 0.1266950, 0.0323755, 0.1057840, 0.0738624, 0.0499694, 0.0696976, 0.0302216, 0.0296763, -0.0406880, -0.0373879, -0.0167024, 0.0024037, 0.0001147, 0.0002060, 0.0015677, 0.0424913, 0.1120170, 0.1913020, 0.2736700, 0.2636380, 0.2116640, 0.3815650, 0.0343093, 0.1581790, 0.1250500, 0.2462350, 0.3790210, 0.2516930, 0.0950500, -0.0311769, -0.0586821, 0.0422582, -0.0341932, 0.1466650, 0.1013130, 0.0979720, -0.0148599, -0.0304525, -0.0061134, 0.0018560, -0.0000581, -0.0007203, -0.0070015, 0.0079964, 0.0655591, 0.1277720, 0.1843750, 0.0688830, -0.0076993, -0.0375187, -0.1282510, -0.0890841, 0.0237801, 0.0881702, 0.1588780, 0.0481340, 0.1611190, -0.0856712, 0.0546686, 0.1963940, 0.1737350, 0.1162280, 0.0213419, 0.0907760, 0.0072640, -0.0132965, -0.0135087, 0.0003164, -0.0001551, -0.0006541, -0.0106625, -0.0230768, -0.0427837, 0.0788373, 0.1291890, -0.0983173, -0.0103092, -0.0494804, -0.0222234, -0.0161273, -0.0589975, 0.1198520, 0.0129883, -0.0454646, 0.2545590, 0.0964659, 0.1759380, 0.0794739, 0.2411300, 0.1061390, 0.0751255, 0.0333420, -0.0205532, -0.0265396, -0.0360304, -0.0000297, -0.0004778, 0.0003995, -0.0039986, -0.0169594, -0.0618618, 0.0050153, 0.1599220, 0.0297676, 0.0202105, -0.0748383, 0.1043680, 0.1473620, 0.1617370, 0.2023150, 0.1251750, -0.0266398, 0.3238990, 0.0758716, 0.1313480, 0.1628160, 0.0641890, 0.0018743, 0.1082160, 0.0854031, 0.0027002, -0.0176384, -0.0290889, -0.0180752, -0.0006609, 0.0003804, -0.0076584, -0.0278685, -0.0197313, 0.0002378, 0.1145280, 0.0755709, -0.0464274, -0.0608713, 0.0132424, 0.0355269, 0.0414473, 0.1112910, 0.0801560, 0.0286425, 0.1180390, -0.0160477, 0.2109670, 0.0272245, -0.0321298, -0.1336420, 0.0601168, 0.0971503, 0.0236622, -0.0685515, -0.0720795, -0.0406126, 0.0001328, 0.0001504, -0.0098816, -0.0271827, -0.0840957, -0.0216471, 0.1034670, 0.1885320, 0.0799817, 0.0878548, 0.1017600, -0.0025078, -0.0366506, 0.3378890, 0.1408050, -0.0231666, 0.1894530, 0.1381170, 0.1199640, 0.1196110, 0.1199460, 0.0507670, 0.1066730, 0.1546050, -0.0908306, -0.1103220, -0.0453135, -0.0081848, -0.0004822, -0.0000498, -0.0032476, -0.0222942, -0.0809317, -0.1083870, 0.0723195, 0.0092438, -0.0978147, 0.1138280, -0.0314414, -0.0234313, 0.0893852, 0.3141660, 0.2549980, -0.0065214, -0.0224469, 0.0408693, 0.0722400, -0.0826778, -0.0228907, 0.0646974, -0.0773966, -0.0543089, -0.1147260, -0.0598585, -0.0183662, 0.0002698, 0.0000206, -0.0000131, -0.0048061, -0.0274983, -0.1290260, -0.1119270, -0.0952378, -0.1091770, 0.0119124, 0.1212930, -0.0683765, 0.1211530, 0.1519980, 0.1228620, 0.0688414, -0.1225560, -0.1233350, -0.2022480, -0.1002740, -0.1211570, -0.0911081, 0.0085364, -0.0331475, -0.0766021, -0.0344098, -0.0406408, -0.0147947, 0.0010590, 0.0002547, 0.0000476, -0.0199242, -0.0720765, -0.0940543, -0.0713264, -0.1638660, -0.1933540, -0.0266128, 0.1817020, -0.0250402, 0.0276831, 0.0466575, -0.1213340, 0.0295884, -0.2678990, -0.2571400, -0.1798960, -0.0139214, 0.0184813, 0.0437714, -0.0602175, -0.0130526, -0.0645854, -0.0270177, -0.0257102, -0.0048713, -0.0000778, -0.0001451, 0.0002514, -0.0324032, -0.0801573, -0.0998883, -0.1191770, -0.2172340, -0.2423570, 0.0103417, -0.0573569, 0.0456261, -0.0432571, -0.1119950, -0.2087320, -0.1091470, -0.0251970, -0.0618544, -0.0294190, 0.0153294, -0.0038500, 0.1203950, -0.0436650, -0.0299444, -0.1076490, -0.0417105, -0.0409794, -0.0071382, -0.0001046, -0.0008609, 0.0002320, -0.0054939, -0.0109514, -0.0030036, -0.0342237, -0.1814830, -0.3181620, -0.2793050, -0.2956670, -0.1193040, -0.0155505, -0.0986209, -0.0683331, 0.0315920, 0.0406260, 0.1212780, 0.0247887, 0.1616530, 0.1226600, 0.0838768, -0.0930329, -0.0564129, -0.0858891, -0.0338816, -0.0426510, -0.0051800, 0.0000304, -0.0000902, 0.0005889, 0.0004757, 0.0234311, -0.0201526, 0.0333871, -0.0928994, -0.1922910, -0.0281642, -0.2837330, -0.2926960, -0.3722260, -0.2181620, 0.0442903, 0.0042594, 0.0298694, 0.0237936, 0.1964730, 0.2590500, 0.1700880, 0.0719090, -0.0589024, -0.0449341, -0.0646688, -0.0359445, -0.0415502, 0.0001586, 0.0004717, 0.0001508, -0.0001930, 0.0012566, 0.0045470, -0.0289076, -0.0728262, -0.1056090, -0.0788080, -0.0183602, -0.1538390, -0.0303134, 0.0387993, -0.1036640, -0.2757910, -0.0919790, -0.0831569, 0.1709660, 0.0921235, 0.0059665, 0.1021750, 0.1225060, 0.0548892, 0.0579596, 0.0426221, -0.0404542, -0.0171239, -0.0020878, 0.0000519, -0.0002600, 0.0003592, 0.0001778, -0.0104153, -0.0572517, -0.0040627, -0.0150223, 0.0104719, 0.0680042, -0.0083080, 0.1219150, 0.0715756, 0.1059160, 0.1796630, 0.1441370, -0.0399740, -0.0718035, -0.0660457, -0.0356566, 0.0943911, 0.1200420, 0.0792530, 0.0315256, 0.0099373, 0.0015349, -0.0012851, -0.0021307, 0.0002662, 0.0004242, 0.0004547, -0.0004520, -0.0002627, 0.0124197, 0.0950441, 0.0908244, 0.0010337, -0.0435880, -0.0571582, -0.0075926, 0.0927066, 0.0811021, -0.0170540, -0.0462112, -0.0888039, -0.0828597, 0.0075775, -0.0320296, -0.0391621, 0.0009601, 0.0048586, -0.0016904, -0.0002353, 0.0006032, -0.0005606, -0.0003848, 0.0007397, -0.0000276, 0.0003083, -0.0001918, -0.0004274, 0.0005511, 0.0002518, -0.0006003, 0.0002914, -0.0002797, -0.0014979, -0.0063987, -0.0029212, -0.0015570, -0.0014733, 0.0051354, 0.0009391, -0.0013568, -0.0004309, 0.0055687, 0.0012160, 0.0008829, 0.0008743, 0.0037383, -0.0006011, -0.0003864, 0.0001110, 0.0001496, 0.0005402, 0.0006172, 0.0001828, 0.0006909, -0.0006454, -0.0003025, 0.0001366, 0.0001978, -0.0000974, 0.0001515, -0.0004436, 0.0004282, -0.0003418, 0.0003571, 0.0006852, -0.0001127, -0.0004795, -0.0002898, 0.0004085, 0.0002279, 0.0004386, -0.0000957, 0.0002139, -0.0000136, 0.0003142, 0.0000652, -0.0006361, 0.0004573, 0.0001703, 0.0002870, 0.0001493, 0.0007542, -0.0000498, -0.0003031, -0.0003050, -0.0002510, 0.0003865, 0.0006532, 0.0015481, 0.0063107, 0.0065363, 0.0047900, 0.0011893, -0.0023838, 0.0032039, -0.0083129, 0.0015414, 0.0039626, 0.0121842, 0.0203436, 0.0091888, 0.0004003, -0.0003247, -0.0000039, -0.0006345, 0.0002581, -0.0004930, 0.0004913, 0.0005550, 0.0002259, 0.0001960, 0.0011444, 0.0005863, 0.0019253, 0.0037659, -0.0008778, -0.0328847, -0.0426598, -0.0092137, -0.0053171, -0.0388914, -0.0455082, -0.0313261, -0.0110661, 0.0329317, 0.0357186, 0.0433980, 0.0318446, 0.0305573, 0.0178815, 0.0073109, -0.0062437, -0.0059448, 0.0000525, -0.0002531, -0.0004907, -0.0005166, -0.0038839, -0.0012675, 0.0037514, -0.0102282, -0.0101183, -0.0141179, -0.0444495, -0.0688281, -0.1498070, -0.2143800, -0.2213880, -0.1466550, -0.0700918, -0.0456266, -0.1020770, -0.0538809, 0.1317900, 0.0771036, 0.0912988, 0.0977176, 0.0705981, 0.0440365, -0.0069990, 0.0017092, 0.0040501, 0.0002943, 0.0004974, -0.0000046, -0.0128910, -0.0051699, -0.0027806, -0.0336706, -0.0195392, 0.0194954, -0.1575900, -0.2018330, -0.2302120, -0.2330970, -0.2501070, -0.1757710, -0.0610809, -0.0550162, -0.0515459, -0.0840172, -0.1276020, 0.0101861, 0.0022437, 0.1145270, 0.0952536, 0.1605650, 0.0607997, 0.0295550, 0.0041381, 0.0026861, -0.0004694, 0.0000946, -0.0045678, -0.0049654, -0.0231581, -0.0436363, -0.0250587, -0.1661450, -0.2016600, -0.1578080, -0.0444237, -0.1593070, -0.2645350, -0.1732470, -0.0822259, -0.0636970, -0.0635151, 0.0173707, -0.1525260, -0.0859735, -0.0638592, -0.0119553, 0.0497776, 0.0705422, 0.0420119, 0.0350166, 0.0097057, 0.0041052, 0.0002225, -0.0001324, -0.0037171, -0.0320082, -0.1179680, -0.1963750, -0.2452970, -0.2602760, -0.0369206, -0.1415290, -0.2336370, -0.3506420, -0.2399480, -0.2995200, -0.1611880, -0.1344780, 0.0144744, -0.0189761, -0.1658860, -0.1026190, -0.1234280, -0.1637440, -0.0446738, 0.0995109, 0.0120174, 0.0341479, 0.0037373, 0.0034115, 0.0000815, -0.0093644, -0.0012191, -0.1154210, -0.2313460, -0.1871660, -0.2644440, -0.2305260, -0.1825160, -0.1864430, -0.0747279, -0.4452160, -0.2977970, -0.3019530, -0.3067320, -0.0034584, -0.1121340, -0.0682714, -0.0473488, 0.0246074, 0.0903544, 0.0848562, 0.0347291, 0.0091155, 0.0573025, 0.0779422, 0.0102823, 0.0012743, 0.0003391, -0.0065070, 0.0077438, -0.0599938, -0.1827400, -0.0686432, 0.1051030, -0.0330234, -0.0340820, -0.1063600, -0.1645840, 0.0375006, -0.0231350, 0.0313613, -0.0583751, -0.0710633, -0.0040034, -0.0403435, 0.0926855, 0.0709464, 0.0426386, 0.1012800, 0.0901951, 0.0779442, 0.1352980, 0.0958148, 0.0096213, 0.0002527, -0.0001765, -0.0030258, -0.0070812, -0.0073654, -0.0770139, 0.1076570, 0.2438870, 0.1105560, 0.2429400, 0.4911130, 0.7808800, 0.8365580, 0.7849860, 0.6271240, 0.1595360, 0.0950786, 0.1724670, 0.1021930, 0.0140080, 0.1500770, 0.0863036, 0.0426656, -0.0167842, -0.0061895, 0.1438350, 0.0194806, 0.0222658, 0.0021590, -0.0005765, -0.0023402, -0.0169275, -0.0136975, 0.1575750, 0.4472910, 0.6555300, 0.9350330, 1.2476500, 1.4381800, 1.1881000, 0.9072770, 0.6861270, 0.3340640, 0.1274250, 0.2727330, -0.0814077, -0.0653220, -0.1242420, 0.0544268, -0.0299599, 0.0127470, 0.0044352, 0.0304259, 0.1016880, 0.0190889, 0.0129452, -0.0012662, 0.0001529, -0.0036237, -0.0719993, -0.0427465, 0.1416630, 0.4904890, 0.6964780, 0.8753270, 0.9015370, 0.6802880, 0.2453460, -0.0438393, -0.1530760, -0.1375150, -0.2091280, 0.0382348, 0.1615570, -0.0009761, 0.0767798, -0.0273172, -0.1202590, 0.1300290, 0.0511068, 0.0401559, 0.0830926, 0.0415490, 0.0217123, -0.0046027, 0.0000496, -0.0010880, -0.0445179, -0.0322498, 0.1424920, 0.2032540, 0.3098000, 0.2034140, -0.0241976, -0.2152100, -0.5068490, -0.3795330, -0.4930990, -0.1278290, -0.2156040, 0.0574476, -0.0263473, 0.1721090, -0.0389348, 0.0033202, 0.0842200, 0.1299820, 0.0718242, 0.1350290, 0.0022822, -0.0918741, -0.0313514, -0.0144558, -0.0000417, 0.0000998, -0.0356313, -0.1110670, -0.0215535, -0.0847103, -0.1644100, -0.3231990, -0.3609730, -0.4179310, -0.5042630, -0.1624360, -0.0859620, -0.0537205, -0.0867637, 0.0671770, 0.1013200, 0.1122180, -0.1710790, -0.0200284, 0.0257647, -0.0009569, 0.1221010, 0.1754290, 0.0964777, -0.0570247, -0.0182045, -0.0002799, -0.0001587, -0.0003883, -0.0128844, -0.1309650, -0.2048420, -0.1681900, -0.2371130, -0.2927470, -0.1749620, 0.0256156, -0.0010701, 0.0442501, -0.0747489, 0.0298914, -0.1581730, -0.0322517, -0.0127613, 0.0204888, -0.0616515, -0.0035494, -0.0668576, -0.0444659, 0.1396700, 0.1216590, 0.1101040, -0.0619533, -0.0489104, 0.0000552, -0.0006518, -0.0013771, -0.0016916, -0.1093740, -0.1800390, -0.2394620, -0.2622780, -0.0061299, 0.3449920, 0.0531424, -0.0035019, 0.0712339, 0.0229197, 0.0037986, 0.0255992, 0.0090434, -0.0138366, 0.2429920, 0.1152700, 0.0465617, 0.0621921, 0.0386113, 0.1795890, 0.0817529, -0.0106259, -0.0202225, -0.0388053, -0.0109606, -0.0005282, -0.0010689, -0.0061135, -0.1005590, -0.2051840, -0.2045090, -0.0797609, 0.0238650, 0.1509500, -0.0808445, 0.0887981, 0.0821237, 0.1824750, 0.0622324, -0.0913239, 0.0670867, 0.0047924, 0.0858643, -0.0949107, 0.0127151, 0.0396182, 0.0507667, 0.0446282, -0.0439240, -0.0140018, -0.0227924, -0.0643085, -0.0251071, 0.0001241, -0.0006743, 0.0013450, -0.1061460, -0.0672064, -0.0258413, 0.0832080, 0.1024140, 0.0543914, 0.1366010, 0.1039870, 0.0005317, 0.1047640, -0.0123072, 0.0337299, 0.0787247, 0.0702442, 0.1762520, -0.0254464, -0.0016614, 0.1678090, -0.0172795, -0.0704116, 0.0025469, -0.0080458, -0.0666274, -0.0435325, 0.0063766, -0.0025316, 0.0005710, -0.0100826, -0.1139590, -0.0050165, 0.0985650, 0.0877037, 0.0755586, -0.0522449, -0.1300860, 0.0208557, 0.1602730, 0.0630176, 0.0416929, 0.0954576, 0.0184258, 0.1159540, -0.0422802, -0.0049141, 0.0203671, 0.0267828, -0.1920140, -0.1878690, -0.0315761, -0.0197203, -0.0751014, -0.0205508, -0.0072401, 0.0001774, -0.0024971, 0.0142187, -0.0918897, 0.0194573, 0.1190020, -0.0624662, -0.0108846, 0.1000310, 0.0570473, -0.0073708, -0.0646952, -0.2018000, -0.2597750, -0.1094160, -0.0399217, -0.0393269, -0.1206560, 0.0092218, -0.0378979, -0.1171660, -0.1891340, -0.1383650, -0.0688766, -0.0222924, -0.0882502, -0.0407872, -0.0021736, -0.0007510, 0.0072174, 0.0245788, -0.0769862, 0.0590626, 0.0330006, 0.0435863, 0.0879408, 0.0196239, -0.0080216, -0.1224920, -0.0045490, -0.0434923, -0.0194296, -0.2593990, -0.1004100, 0.0111438, 0.0132768, -0.1764110, 0.0212538, 0.0178922, -0.1323280, -0.1087620, -0.0119571, -0.0021344, -0.0337255, -0.0143575, 0.0000834, -0.0001112, -0.0007536, -0.0111720, -0.0323503, 0.0340453, 0.0810478, 0.0159146, 0.0199603, 0.0525500, 0.1672580, -0.0160685, 0.0603623, 0.0872160, 0.1010330, -0.0019192, 0.0463692, -0.1605190, -0.0385112, -0.0435163, 0.0380387, 0.1181280, 0.0688014, 0.0041884, -0.0536306, -0.0389279, -0.0180200, -0.0030185, -0.0004880, 0.0006847, 0.0002440, -0.0074172, 0.0128627, -0.0616254, -0.0748103, 0.0022474, -0.0797940, 0.0506937, 0.0752191, -0.0905753, 0.0280538, 0.0929923, 0.0412421, -0.0571475, -0.0360529, -0.0386100, 0.1216370, 0.1134240, -0.0156331, 0.0128100, 0.1223960, 0.0771567, -0.0040338, -0.0094860, 0.0007675, 0.0005320, -0.0000633, 0.0001391, -0.0007719, -0.0077499, -0.0471869, -0.0624455, -0.0854893, 0.0658057, -0.0508412, 0.0121698, -0.0475049, 0.0838423, -0.0407969, 0.0365388, -0.0609659, 0.0499621, -0.0190625, -0.0515456, 0.0970983, 0.1701280, 0.1072720, 0.1312520, 0.0858693, 0.0146668, -0.0342011, 0.0015156, 0.0030614, -0.0044381, -0.0000601, 0.0002727, 0.0003907, -0.0034983, -0.0464869, -0.0628340, -0.0190867, -0.0990476, -0.1369510, -0.1063720, 0.0029366, -0.0357361, -0.1383710, 0.0841809, 0.0358197, -0.1193890, 0.0678497, 0.0969432, -0.1407190, -0.0072907, 0.0752326, 0.0562790, -0.0506607, -0.0498293, 0.0201849, 0.0001848, -0.0004099, -0.0001699, -0.0004160, 0.0001663, -0.0003112, -0.0006859, 0.0013088, -0.0505133, -0.0532395, -0.0846707, -0.0629257, -0.0794203, -0.0652940, -0.0237631, 0.0152936, -0.0815658, -0.1531030, -0.0450743, 0.1556580, -0.0176126, -0.1644610, -0.1086080, -0.0484371, -0.0138990, 0.0162404, -0.0176824, 0.0082222, -0.0004382, 0.0006892, 0.0012003, -0.0002040, -0.0000155, 0.0003468, 0.0001048, 0.0001551, -0.0045516, -0.0140714, -0.0084642, 0.0252005, -0.0199096, -0.0585476, -0.0843062, -0.0207266, -0.0086491, -0.0454075, 0.0393739, 0.0373841, -0.0722731, -0.0977680, -0.0593750, -0.0495706, -0.0349817, 0.0121983, -0.0060897, 0.0002496, -0.0002147, -0.0000837, 0.0003760, 0.0004731, 0.0002229, -0.0003291, -0.0005079, -0.0002090, -0.0002073, -0.0000265, 0.0010788, 0.0020959, 0.0021280, 0.0011776, 0.0067339, 0.0052072, 0.0014372, 0.0021502, 0.0069564, 0.0004217, -0.0268756, -0.0079765, 0.0025296, -0.0008624, -0.0007181, -0.0000295, -0.0005459, -0.0003488, 0.0002264, 0.0001438, 0.0003744, 0.0005680, -0.0001344, 0.0005911, 0.0000542, 0.0000842, 0.0000235, -0.0000232, 0.0001352, -0.0002237, -0.0003237, -0.0002169, -0.0006377, -0.0000732, 0.0007089, 0.0014808, 0.0001340, -0.0000591, 0.0004927, 0.0004254, -0.0001390, -0.0000946, 0.0001155, 0.0002288, -0.0004770, 0.0002559, -0.0002473, 0.0003599, 0.0002979, 0.0002084, -0.0000138, 0.0008709, 0.0000652, -0.0005757, -0.0007766, 0.0002176, 0.0017550, 0.0031662, 0.0071776, 0.0018322, 0.0057806, 0.0003126, 0.0011888, 0.0005921, -0.0089246, -0.0103576, -0.0210814, -0.0005413, 0.0098279, 0.0101048, 0.0144327, 0.0139610, 0.0014194, 0.0003562, -0.0000366, 0.0003310, 0.0000257, -0.0004972, 0.0004097, -0.0002192, -0.0000377, -0.0002837, -0.0004327, -0.0000217, 0.0030170, 0.0110022, 0.0126570, 0.0049200, 0.0053618, -0.0002061, 0.0096291, -0.0130107, -0.0224744, -0.0364781, -0.0400377, 0.0165447, 0.0151119, 0.0202901, 0.0134911, 0.0254354, 0.0266348, 0.0082172, -0.0008748, -0.0029168, 0.0000678, 0.0000553, -0.0003298, -0.0001856, -0.0043661, -0.0008691, -0.0016510, 0.0003859, 0.0052277, 0.0013909, -0.0477495, -0.0329655, 0.0000532, -0.0574863, -0.1025240, -0.1131880, -0.0668807, -0.0317981, -0.1105600, -0.0973283, -0.0582066, -0.0326379, 0.0471968, 0.0435064, 0.0581568, 0.0453528, 0.0145650, 0.0026276, 0.0072023, 0.0007469, -0.0001786, 0.0000972, -0.0152521, -0.0032596, 0.0046816, -0.0080989, -0.0186801, 0.0023747, 0.0118625, 0.0935688, 0.0839001, 0.0176852, 0.1056810, 0.1176030, 0.1585170, 0.0734982, -0.0302766, 0.0934747, -0.0696782, -0.1525870, -0.1342000, 0.0817646, 0.0488843, 0.0608986, 0.0649226, 0.0205462, 0.0137191, 0.0129645, 0.0003091, 0.0001621, -0.0020357, -0.0053096, -0.0267670, -0.0458394, 0.0103151, -0.0278687, -0.0090464, -0.0898265, -0.0173192, 0.0912187, 0.1005910, 0.0639935, 0.0604582, 0.1059900, -0.1901400, 0.1537530, 0.1000360, 0.0511407, 0.0125859, 0.1168220, 0.0865553, 0.0941551, 0.1090200, 0.0947396, 0.0521279, 0.0191149, 0.0000718, -0.0002024, -0.0020995, -0.0496479, -0.0638129, -0.0914783, -0.1601430, -0.0752998, -0.0111032, -0.1563040, -0.2312110, 0.0712229, 0.1486050, 0.0021598, -0.0850318, -0.0902836, -0.1060660, 0.1382370, -0.0528104, -0.0138788, 0.0982434, 0.2338400, 0.1115420, 0.1815960, 0.1010400, 0.1095660, 0.0283575, 0.0158814, -0.0000646, -0.0107149, -0.0115374, -0.0614539, -0.0627877, -0.0676763, -0.1381380, -0.1400550, -0.0509202, -0.1277050, -0.1689160, -0.1199860, -0.0469921, -0.0890481, -0.0974893, -0.0387921, -0.0643921, -0.1349720, 0.0612303, -0.2681570, -0.1912520, 0.1381770, 0.0326493, 0.1111610, 0.1027980, 0.1153090, 0.0295050, 0.0102316, -0.0002810, -0.0037804, -0.0060930, -0.0249363, -0.0874373, -0.1084050, 0.0129296, -0.1472930, -0.1220560, -0.0401549, -0.1922570, -0.2038880, 0.0675108, -0.0036416, -0.2198100, -0.1170380, 0.0512611, -0.2849990, -0.0746176, -0.0210022, -0.0240782, 0.1400490, -0.0741726, 0.0718466, 0.2507950, 0.1036680, 0.0160487, 0.0013007, 0.0001831, -0.0029937, -0.0125299, -0.0163207, -0.0516998, -0.1444410, -0.0645730, -0.2498200, -0.2769860, -0.2051910, -0.2083240, -0.1731580, -0.2575460, 0.1614410, 0.1111590, -0.1021910, -0.0564832, 0.0013058, 0.0423332, 0.1966350, 0.2624340, 0.1235750, -0.1523640, 0.1249370, 0.1976050, 0.0851070, -0.0212696, -0.0539882, 0.0001334, -0.0014968, -0.0029367, 0.0053111, 0.0783083, 0.0281975, -0.0217701, -0.2823250, -0.3394460, -0.0548348, -0.1058220, 0.0798663, 0.3597790, 0.5137420, 0.6317750, 0.1424530, -0.1219030, -0.0568714, -0.0200343, 0.0723104, 0.0934951, 0.0527661, 0.1556220, 0.1439470, 0.0687969, -0.0469861, -0.0297524, -0.0165617, 0.0002226, -0.0004680, 0.0209829, 0.0489655, 0.2350720, 0.2614850, 0.2183170, 0.2799040, 0.3018220, 0.6307560, 0.8020010, 0.9173870, 1.3766000, 0.9182140, 0.4178720, 0.0517402, -0.0650657, -0.0207738, 0.0622322, -0.0502315, -0.0375738, 0.0410937, 0.1027190, 0.1689010, 0.1166690, -0.0169929, 0.0404969, 0.0006702, 0.0002181, 0.0008324, 0.0121284, 0.0943970, 0.3409860, 0.4808890, 0.5987820, 0.8587670, 1.0741900, 1.4377100, 1.0918100, 0.9390710, 0.4769650, 0.1288290, 0.0591672, 0.0139135, -0.1108840, 0.0221528, -0.0183021, 0.1538440, 0.0273881, 0.1011360, 0.1712540, 0.2131140, 0.1524670, -0.1257080, -0.0181563, -0.0037547, 0.0006260, 0.0010231, -0.0045445, 0.1088060, 0.4000380, 0.7906600, 0.8031860, 0.9664390, 0.9095280, 0.6788640, 0.3698300, 0.1118970, -0.1856640, -0.1576200, -0.0143233, 0.0586130, 0.0239192, 0.0267489, 0.0925160, 0.1603440, 0.1736220, -0.0211592, 0.0468735, 0.0308513, -0.0796043, -0.1875970, -0.0630238, -0.0159337, -0.0002782, -0.0022499, -0.0082612, 0.1047680, 0.2661720, 0.5531720, 0.4212450, 0.3405330, 0.2202840, -0.1983190, -0.3614060, -0.2877330, -0.3807320, -0.2079110, -0.2528950, -0.1573650, -0.0736923, -0.0415607, -0.1333550, -0.0523307, -0.0081361, -0.0699596, -0.0550363, -0.1767730, -0.1793830, -0.1337680, -0.0674149, -0.0019257, -0.0005340, -0.0045565, -0.0041471, 0.0232957, 0.1167730, 0.1430210, 0.0354759, -0.1556640, -0.2073610, -0.1371080, -0.1532870, -0.0619865, -0.1010020, -0.2027840, -0.0980110, -0.1516870, 0.0193071, 0.0001051, -0.2299250, -0.0287865, 0.0273164, -0.1664460, -0.0429344, -0.1759220, -0.1507160, -0.0417561, -0.0115251, -0.0032804, -0.0003340, -0.0029096, -0.0147998, -0.0919453, -0.0251999, -0.0587297, -0.1663140, -0.2559260, -0.1045800, 0.0200354, -0.0186940, -0.0412775, -0.0769017, -0.1858630, -0.0575565, 0.0368003, 0.0105433, 0.0269425, -0.1625770, -0.2738050, -0.0633486, -0.1327580, -0.0493528, -0.1479870, -0.2251130, -0.0561205, -0.0565053, -0.0085663, -0.0005101, -0.0002075, -0.0169033, -0.1288060, -0.1763390, -0.0902387, -0.1209160, 0.0192422, 0.0611677, 0.0144881, 0.0287163, 0.0075700, -0.2045120, -0.1824210, -0.1509420, -0.0758979, -0.0059501, 0.0557734, -0.0089214, -0.1711770, 0.1461110, 0.0049938, -0.0373651, -0.0471809, -0.0769919, -0.0464294, -0.0418005, -0.0122991, -0.0002541, -0.0001715, -0.0119529, -0.1545770, -0.1742080, -0.1327080, -0.0713065, 0.0466169, 0.0454337, -0.0760951, -0.0340469, -0.0506673, -0.2327090, -0.0653244, -0.1106420, -0.1414550, -0.0772552, -0.1137920, -0.0046588, -0.0942593, 0.1573710, 0.1239310, 0.0542168, 0.0392663, -0.0807243, -0.1163260, -0.0282723, -0.0116214, -0.0001005, 0.0026393, -0.0052296, -0.0573370, -0.1783390, -0.0856638, -0.2007410, -0.1578330, 0.0665130, -0.0172350, -0.0512633, -0.0986202, 0.0324762, -0.1204160, 0.0481937, 0.0343921, 0.0033982, -0.0975658, 0.1477920, 0.0407908, 0.0811889, -0.0547952, 0.0383914, 0.0477377, -0.0386766, -0.1048640, -0.0059238, -0.0029222, -0.0005586, 0.0075830, -0.0092031, -0.1520500, -0.1727590, -0.1652550, -0.1631200, -0.0197090, 0.0279196, -0.0787290, 0.0353450, -0.0356574, 0.0859175, 0.0898348, -0.0946055, 0.0328007, 0.0325335, 0.0296671, 0.0109885, -0.0693787, -0.0362466, -0.0561792, 0.0948938, 0.0732430, 0.0062063, -0.0666466, -0.0038788, 0.0002924, -0.0003079, -0.0004446, -0.0255462, -0.1515050, -0.0767313, -0.1170160, 0.0250049, -0.0440897, 0.0146693, 0.0168059, -0.0984152, 0.0161136, -0.1589070, -0.0937304, -0.0406523, -0.0583694, -0.0129666, -0.0054170, -0.0723663, -0.1071730, 0.0482405, -0.0679664, 0.1446170, 0.0806481, -0.0290826, -0.0443066, -0.0024626, -0.0003275, 0.0004654, 0.0000750, -0.0223371, -0.0307185, -0.1634950, -0.2350060, 0.0762570, -0.0502542, -0.0787612, 0.0934066, 0.0755301, 0.0021196, 0.2231520, -0.0740215, -0.0392414, -0.0351312, -0.2291160, -0.0135183, 0.0569305, -0.1052800, -0.0357939, 0.0523001, 0.1484900, 0.0701413, -0.0124337, -0.0250431, -0.0047780, 0.0005792, 0.0002231, 0.0002354, -0.0033266, -0.0199932, -0.1081600, -0.2657220, -0.1783670, -0.1935610, -0.0305720, -0.0454785, 0.2454320, 0.0290295, -0.0006737, -0.1712620, 0.0811819, -0.0522163, -0.0058234, 0.0743493, -0.0060774, 0.0345833, 0.0726968, 0.0645144, 0.0795196, 0.0471677, -0.0259689, -0.0212113, -0.0048576, 0.0001928, 0.0001549, -0.0001512, -0.0005818, -0.0234185, -0.0923864, -0.1074460, 0.0052725, 0.0135535, -0.0426803, -0.0871856, 0.0332209, 0.0280994, 0.0616517, 0.1579350, 0.0711563, 0.1077160, 0.1530820, -0.0759414, 0.1677900, 0.2008490, 0.0443109, 0.0520710, 0.0512092, 0.0204015, -0.0516615, -0.0076851, -0.0029556, 0.0000888, 0.0000235, -0.0005669, 0.0007268, -0.0154824, -0.0469201, 0.0196229, -0.0047692, -0.0441377, -0.1050850, -0.0748203, -0.0632865, -0.0122861, -0.0807010, 0.1778650, 0.0464078, -0.1588350, -0.0896681, 0.0468261, 0.2019790, 0.1323980, 0.0507034, 0.1152520, 0.0624963, 0.0164736, -0.0005854, -0.0027307, -0.0023415, 0.0000666, -0.0004290, 0.0003125, 0.0004888, -0.0001483, 0.0210681, 0.1411320, 0.1221030, -0.0045150, -0.0181719, -0.0218804, -0.0237605, 0.0001142, 0.0268807, 0.0284220, -0.0179389, -0.0091602, 0.0607794, 0.0221002, -0.0037227, 0.0068307, 0.0205543, 0.0607540, 0.0336342, 0.0005137, -0.0001485, -0.0001648, 0.0001729, 0.0000017, 0.0002427, -0.0000905, -0.0003739, -0.0001589, -0.0007151, -0.0004059, -0.0007669, -0.0006538, -0.0010591, -0.0035456, -0.0123428, -0.0055191, -0.0021712, -0.0016435, 0.0004761, -0.0022105, -0.0018090, -0.0104297, -0.0126396, 0.0053567, 0.0064457, 0.0061150, 0.0403480, -0.0005505, -0.0001592, 0.0002989, -0.0001292, 0.0001080, -0.0000211, -0.0001760, 0.0000045, 0.0000791, -0.0000217, 0.0000864, -0.0003225, 0.0007898, 0.0002898, -0.0001447, 0.0003560, 0.0007326, 0.0010959, 0.0033454, -0.0006192, 0.0001060, 0.0000147, 0.0001193, -0.0001156, -0.0005475, 0.0000623, -0.0004862, -0.0002188, -0.0003482, 0.0006598, -0.0003636, -0.0002654, -0.0002678, -0.0000871, 0.0000177, 0.0001895, -0.0004898, 0.0003778, 0.0005979, 0.0004517, 0.0004770, -0.0011813, -0.0009654, -0.0008750, 0.0005485, 0.0027979, 0.0000892, 0.0046793, 0.0016739, -0.0142707, -0.0056722, -0.0003833, 0.0002958, 0.0007974, 0.0014017, 0.0002139, -0.0001290, 0.0000408, -0.0004391, -0.0004506, -0.0004255, -0.0002944, -0.0000295, 0.0002407, -0.0014010, -0.0007523, -0.0001727, 0.0020213, 0.0028292, 0.0055088, 0.0274183, 0.0128680, 0.0225213, 0.0264469, 0.0461351, 0.0667633, 0.0537765, -0.0037635, -0.0088322, -0.0094574, -0.0061461, -0.0079506, 0.0044022, 0.0035216, -0.0049112, -0.0043852, -0.0027371, 0.0004782, -0.0001973, 0.0000142, -0.0000841, 0.0000679, -0.0048879, -0.0008147, 0.0049217, 0.0063094, 0.0176704, 0.0188385, 0.0416864, 0.0405001, 0.0514171, 0.0211103, 0.0746670, 0.1798670, 0.1281970, 0.0563606, -0.0009563, -0.0184586, 0.0291454, 0.0093178, 0.0066226, -0.0006775, -0.0095680, -0.0068001, -0.0020218, 0.0001087, 0.0001628, -0.0002319, 0.0000313, -0.0005997, -0.0006028, 0.0025992, 0.0251287, 0.0295988, 0.0769531, 0.1465370, 0.1439080, 0.1728320, 0.0958467, 0.0940411, 0.2111720, 0.1436100, 0.0720360, 0.1065550, 0.0408681, -0.0058425, 0.0057574, 0.0029575, 0.0028644, 0.0382182, -0.0182298, -0.0376771, -0.0113300, 0.0089661, 0.0083246, 0.0005314, -0.0005068, -0.0001713, -0.0007288, 0.0127978, 0.0230878, 0.0731718, 0.1639050, 0.2202860, 0.2073450, 0.2604200, 0.0732613, 0.3554040, 0.4839310, 0.5985420, 0.3964460, 0.2843340, 0.3287080, 0.1582890, 0.1589940, 0.1105520, 0.0896389, 0.1265100, 0.1072340, 0.0808457, 0.0807332, 0.0262778, 0.0124986, 0.0003910, -0.0004637, -0.0004988, -0.0604423, -0.0537323, 0.0064226, -0.0121213, 0.1011250, 0.1908020, 0.1761860, 0.1579760, 0.0901179, 0.2321980, 0.0724445, 0.3475470, 0.6455820, 0.6793210, 0.4910600, 0.5307350, 0.4131610, 0.4235530, 0.2114860, 0.2030530, 0.1926090, 0.1221890, 0.0941684, -0.0101805, -0.0030451, -0.0000600, -0.0004068, -0.0011627, -0.0767085, -0.0452845, 0.0502267, -0.1213240, -0.1069810, -0.1429900, 0.0152084, -0.0998191, -0.0246290, -0.0637299, -0.1351230, 0.0579613, 0.2464980, 0.5391560, 0.6555180, 0.7460740, 0.5334190, 0.2933300, 0.1848370, 0.0786049, 0.0512362, 0.0123054, 0.0303885, -0.0018439, -0.0024228, 0.0012331, -0.0017346, 0.0003233, -0.0222973, -0.0224366, 0.0135828, -0.1071680, -0.0404498, -0.0598643, -0.0116079, -0.3656050, -0.1827680, -0.1351040, -0.1127880, 0.0311304, -0.0375656, 0.1339060, 0.0460941, 0.1453270, -0.0759121, -0.0687449, -0.0325362, -0.0141339, -0.1272190, -0.2018220, -0.0097557, -0.0227594, -0.0059536, 0.0003436, -0.0021008, -0.0016303, -0.0211087, -0.0661305, -0.0704463, -0.1995730, -0.2212210, 0.0124478, -0.1662600, -0.2040060, -0.1779860, -0.1851940, -0.2890140, -0.3710510, -0.3696660, -0.3950570, -0.5002660, -0.2297520, -0.0918611, 0.1073370, 0.0822183, -0.0744997, -0.0684594, -0.1758780, -0.1024870, -0.0851800, -0.0269717, -0.0000552, -0.0012477, -0.0042761, -0.0489021, -0.0679073, -0.1072360, -0.3712410, -0.0879425, 0.0695933, -0.1620710, -0.1742100, -0.1342280, -0.1058360, -0.4152340, -0.4719190, -0.3808510, -0.6334620, -0.2640040, 0.0035965, -0.0079745, -0.0247578, 0.0938159, -0.0497112, -0.0877583, -0.0888940, -0.1613760, -0.0722597, -0.0079618, -0.0002467, -0.0018791, -0.0509525, -0.0954186, -0.1530110, -0.1311370, -0.2129580, -0.0187425, -0.0187185, -0.1080860, -0.0265863, -0.3090910, -0.1896600, -0.3363600, -0.2659570, -0.3642720, -0.3237170, -0.2590790, -0.0693696, -0.1135440, -0.0835543, 0.0478209, -0.1243280, -0.0023894, -0.1233670, -0.0935000, -0.0291922, -0.0043723, -0.0000543, -0.0012138, -0.0199139, -0.0901319, -0.1882350, -0.0559372, -0.0624456, -0.1772620, -0.1519330, -0.1072060, 0.2114370, -0.0347356, 0.1516690, -0.0602641, -0.1910010, -0.1127860, -0.0265405, -0.2604760, 0.1385700, 0.0904100, 0.1727500, 0.1207570, 0.0883171, 0.1620550, 0.1129440, -0.0926181, -0.0832077, -0.0123668, 0.0002241, -0.0007343, -0.0135692, -0.0597816, -0.1202050, 0.0374222, -0.0436939, -0.0155919, 0.1614680, 0.2059220, 0.2628690, 0.0172278, 0.1376630, 0.1434970, 0.1718540, 0.1902050, -0.0323444, 0.0262964, 0.2368350, 0.2791370, 0.0125164, 0.0244068, 0.0786315, 0.1520870, 0.0020132, -0.1032250, -0.0829409, -0.0070383, 0.0003878, -0.0005058, -0.0046482, -0.0260720, -0.0124019, 0.2608930, 0.0538375, 0.1590720, 0.1267940, 0.0191608, 0.2168270, 0.0656536, 0.1149800, 0.1843490, 0.3300960, 0.1568910, 0.1165360, 0.0919979, -0.0018571, 0.2582140, 0.0446383, 0.1103080, 0.0768020, -0.0040731, -0.1228450, -0.0837761, -0.0540042, -0.0010366, -0.0004497, 0.0003916, -0.0004674, 0.0234998, 0.0008347, 0.0502948, -0.0052746, 0.1432330, -0.0316681, -0.1000540, 0.0070028, -0.0724110, -0.0027590, 0.2002100, 0.1875680, 0.1915450, 0.1402320, -0.0682058, -0.0568475, 0.0022560, 0.0468309, -0.0284916, 0.1494750, -0.0430610, -0.1793090, -0.0414960, 0.0399245, -0.0073234, 0.0002717, 0.0009736, -0.0004786, 0.0088173, -0.0422298, -0.0280212, 0.0371854, -0.0053603, -0.0224157, 0.0242387, 0.0128540, -0.0063779, 0.0145299, 0.1061420, 0.2208790, 0.2729760, 0.2036380, 0.2360830, 0.1123990, -0.0640421, 0.0442862, -0.0087222, -0.0554244, -0.1188360, -0.0414230, 0.0238158, -0.0418885, -0.0192921, -0.0003079, -0.0000894, -0.0008150, -0.0106196, 0.0170309, -0.0601430, -0.0805238, -0.0083055, -0.0097117, 0.0619651, -0.0012279, -0.0192167, -0.1657120, 0.0614465, 0.0903403, 0.0112430, 0.1599420, 0.1324200, 0.0697163, -0.0896089, -0.0271154, 0.0433166, -0.0457295, -0.0708919, -0.0488445, 0.0516015, -0.0122985, -0.0070931, -0.0009647, -0.0001158, -0.0026754, 0.0260105, 0.0779597, -0.1253980, -0.1367930, -0.0134732, -0.0852821, 0.0979257, 0.0400102, -0.1626040, -0.0152574, 0.1095040, 0.0881855, 0.0338351, 0.1413840, 0.0507490, 0.0794237, 0.0249250, 0.0841233, 0.0637082, -0.1364100, -0.0552496, -0.0390479, 0.0035680, -0.0063923, -0.0000422, 0.0004481, -0.0145038, -0.0035018, 0.0386092, 0.0056404, -0.0972382, -0.1187920, -0.1593430, -0.0128829, 0.1324260, 0.0961500, 0.0509897, 0.0268070, 0.1404280, -0.0680444, 0.0713436, 0.0253552, -0.0584507, -0.0200253, -0.0228259, 0.0824211, 0.0056246, -0.0265455, -0.0296683, -0.0587449, -0.0237326, -0.0024826, 0.0001201, 0.0000747, -0.0002280, 0.0007384, 0.0028643, -0.0382462, -0.1230520, -0.1088650, -0.0610999, -0.1810630, -0.0408520, -0.0168030, 0.1581850, 0.2408000, 0.1439650, 0.2380700, 0.2648820, 0.1216580, 0.0998664, 0.0341723, -0.0188637, 0.0521695, 0.0414300, 0.0757346, -0.0587621, -0.0659174, -0.0437108, -0.0001600, 0.0001667, 0.0005298, 0.0004769, 0.0022613, 0.0150188, -0.0284734, -0.0568057, 0.0026748, 0.1520090, 0.0945692, -0.0301520, 0.1070800, 0.1850810, 0.1705800, 0.2439660, 0.3571790, 0.1666920, 0.2267290, 0.2823100, -0.0146420, 0.0323666, 0.0684995, 0.0052152, 0.0392603, -0.0299875, -0.0375055, -0.0459020, 0.0002726, -0.0005202, 0.0005514, -0.0002826, 0.0009685, 0.0022114, 0.0087252, 0.0498635, 0.0830668, 0.1866780, 0.1859840, 0.0076321, 0.1583500, 0.2067090, 0.0365822, 0.0435188, -0.0167997, 0.0550143, 0.1415720, 0.0802768, -0.0518248, 0.2355770, -0.0653472, -0.0298479, -0.0060532, -0.0057778, -0.0317078, -0.0264237, 0.0016271, 0.0000475, -0.0001267, 0.0001735, 0.0006001, -0.0050267, 0.0182143, 0.0256858, 0.1093600, 0.1571840, 0.1701460, 0.2219630, 0.1578290, -0.0233359, -0.0187320, -0.0768506, -0.1366230, -0.1639910, -0.1388640, 0.0266861, 0.1496500, 0.2702130, 0.0068499, 0.0506629, 0.0207279, 0.0225818, 0.0040245, -0.0004676, 0.0005012, 0.0000789, 0.0000819, 0.0002673, 0.0001868, -0.0012479, 0.0017633, 0.0129059, 0.0406416, 0.1018010, 0.1775360, 0.2616580, 0.0549462, 0.0945832, 0.1643000, 0.1722550, 0.1322750, -0.0844416, 0.0220475, -0.0576307, 0.1536150, 0.0897974, -0.0883452, 0.0268841, -0.0160478, -0.0396386, -0.0159098, 0.0029036, 0.0011739, -0.0010053, -0.0001870, 0.0001409, 0.0000472, -0.0012535, 0.0032293, -0.0066943, -0.0438939, -0.0439954, 0.0458640, 0.1342270, 0.0136249, 0.0795158, 0.0035993, -0.0167530, -0.1310760, -0.1312400, -0.2215670, -0.2537060, -0.1563850, -0.2663720, -0.1564370, -0.0982204, -0.0296622, 0.0183037, -0.0045321, 0.0007935, 0.0007045, 0.0001137, 0.0000625, 0.0002914, -0.0003946, -0.0000850, 0.0042948, -0.0081110, -0.0341615, -0.0417540, -0.0267097, -0.0265531, -0.0459858, -0.0962676, -0.1414300, -0.1968090, -0.1615140, -0.1041380, -0.1623020, -0.1613310, -0.1672120, -0.1798400, -0.1120070, -0.0456028, -0.0074607, -0.0013639, -0.0001096, 0.0004020, 0.0002123, 0.0001830, 0.0004645, -0.0003944, -0.0002929, -0.0000886, 0.0002842, 0.0006724, -0.0030248, -0.0209261, -0.0186838, -0.0033188, -0.0172633, -0.0076766, -0.0036314, -0.0053980, -0.0383227, -0.0042036, -0.0286703, -0.0146284, -0.0193760, -0.0044323, -0.0003020, -0.0019407, -0.0023012, -0.0002460, 0.0000243, 0.0000396, -0.0004755, -0.0001108, -0.0001865, -0.0000963, 0.0005625, 0.0003946, 0.0006956, 0.0003639, 0.0006567, -0.0000276, -0.0004520, -0.0000669, 0.0000037, -0.0000975, 0.0007030, 0.0014376, -0.0005892, -0.0002769, 0.0003324, -0.0004713, 0.0001761, 0.0000189, 0.0002990, -0.0004112, -0.0001506, 0.0000431, -0.0004465, 0.0004114, 0.0002805, -0.0000531, -0.0000060, -0.0003909, -0.0000924, -0.0000269, 0.0000322, 0.0002080, 0.0009494, 0.0015838, 0.0022254, 0.0013457, 0.0010934, 0.0003603, 0.0017170, 0.0030382, 0.0124075, 0.0247544, 0.0117874, 0.0146017, 0.0118920, 0.0083881, 0.0120240, 0.0058655, 0.0044703, 0.0001047, 0.0001032, -0.0000988, 0.0001679, 0.0000439, -0.0000893, 0.0011542, -0.0008577, -0.0006571, 0.0006657, 0.0002127, 0.0031390, 0.0068134, 0.0059209, -0.0146673, -0.0355035, -0.0123145, -0.0332558, -0.0440808, -0.0458630, 0.0085131, -0.0111234, -0.0298962, -0.0202113, 0.0327270, -0.0065963, -0.0101764, 0.0021585, 0.0004347, -0.0016239, -0.0003441, -0.0001774, 0.0001014, -0.0001565, 0.0004124, -0.0022906, -0.0003313, 0.0029296, 0.0007119, 0.0060323, 0.0031102, -0.0074944, -0.0087019, -0.0289320, -0.1069550, -0.1239030, -0.2322800, -0.2155240, -0.1126890, -0.0970015, -0.0640258, -0.1560500, -0.0499299, -0.0727624, -0.0566642, -0.0429774, -0.0297228, -0.0117868, 0.0030893, 0.0013275, 0.0003984, 0.0002259, 0.0001070, -0.0082696, -0.0018600, 0.0030651, -0.0011772, -0.0479977, -0.1000690, -0.0631505, 0.0028811, 0.0424039, -0.0230351, -0.0937734, -0.0914754, -0.2696430, -0.2189340, -0.1986360, 0.0225553, -0.0057861, -0.0023943, 0.0154204, 0.0157257, -0.0398071, 0.0893058, 0.0034106, 0.0003440, -0.0025500, -0.0009490, 0.0000231, 0.0000706, -0.0022203, -0.0016291, 0.0127313, 0.0048297, -0.0133460, -0.0413031, 0.0678707, 0.1297180, 0.2835210, 0.2989030, 0.1918390, 0.0860399, -0.0685800, -0.1612430, -0.1265340, 0.0238319, -0.0754409, -0.2703140, -0.2006200, -0.0642890, -0.0277895, 0.1081380, 0.0167231, -0.0177579, -0.0079460, -0.0002712, -0.0002788, -0.0002746, 0.0022715, -0.0172255, 0.0016792, 0.0285083, 0.0541473, 0.0905496, 0.0867971, 0.0509246, 0.0935058, 0.2274070, 0.2222160, 0.0462878, 0.1424030, -0.1374930, -0.1025260, 0.0749857, -0.0281006, -0.2417560, 0.0585949, -0.1056760, -0.1008190, -0.0239695, 0.0087286, -0.0094041, 0.0071064, -0.0000471, -0.0005911, -0.0090404, 0.0038417, -0.0272198, -0.0465462, 0.0190530, -0.0342824, -0.0904384, -0.1111990, -0.0873643, -0.0765856, 0.0200936, 0.0540862, 0.0706867, 0.1748870, 0.0133564, 0.1796920, 0.1176150, -0.1067720, -0.2336010, 0.0339861, -0.0772245, -0.0081576, 0.0555059, 0.0279559, -0.0178750, -0.0052142, -0.0000179, 0.0010166, -0.0019771, 0.0101730, -0.0113042, -0.0863361, -0.0009572, -0.1215450, -0.1242820, -0.0292083, -0.2759400, -0.2917430, -0.2399810, -0.1380130, 0.1129490, 0.2735670, -0.0175490, 0.0333524, -0.2300550, -0.2424640, -0.3094830, -0.0314601, -0.0246729, -0.0885667, -0.0482349, 0.1099390, 0.0152962, -0.0265497, -0.0023698, -0.0000026, -0.0007090, 0.0044015, -0.0328926, -0.0769254, -0.0450809, -0.1045810, -0.1268760, -0.1351680, -0.1389920, -0.0795261, -0.1431930, -0.1492700, 0.1392970, 0.2669590, 0.0812191, 0.0275525, -0.1955840, -0.0404431, -0.0666016, -0.0102835, -0.0689024, -0.2122230, -0.0670599, 0.0842078, 0.0206328, -0.0247128, 0.0027311, 0.0002952, -0.0006232, 0.0067664, -0.0218138, 0.0350900, -0.0808363, -0.1102540, -0.1194150, -0.0002467, 0.0973886, 0.0386242, -0.0051932, 0.3427370, 0.2515680, -0.2001270, -0.0832655, 0.0386065, -0.0631542, -0.1208320, -0.2085030, -0.1280960, -0.1990800, -0.2337030, -0.0283875, 0.1071000, 0.0319935, -0.0357478, -0.0062651, 0.0005391, 0.0006230, 0.0077447, 0.0069793, 0.0845137, 0.1048480, 0.1167310, -0.0137057, 0.0881270, 0.1605380, 0.2417520, 0.3663590, 0.4051560, -0.1532730, -0.6404640, -0.2720430, 0.2084890, 0.1240280, -0.0399440, -0.1610770, -0.1440020, -0.1167030, -0.1174400, -0.0067781, -0.0662822, -0.0809036, -0.0447363, -0.0052170, 0.0003076, 0.0009032, 0.0060525, 0.0531066, 0.1941890, 0.3282070, 0.3921770, 0.2907770, 0.3347770, 0.3355510, 0.2703880, 0.1426900, -0.0635876, -0.4282140, -0.4729640, -0.0862561, 0.1520520, -0.0053859, 0.1462960, 0.0152932, -0.0766193, -0.0778089, 0.0960453, 0.1099140, -0.0792374, -0.1039860, -0.0424148, -0.0044330, 0.0004035, 0.0019381, -0.0007042, 0.0098972, 0.2319610, 0.3722920, 0.4520510, 0.5285410, 0.2005420, 0.2346810, 0.3065910, -0.0790222, -0.2010570, -0.3632140, -0.0414229, 0.0885448, -0.0998328, -0.0441672, 0.1817170, 0.0722460, -0.0888804, 0.1388590, 0.1305140, 0.1281010, -0.0626949, -0.0897707, -0.0683660, -0.0116694, 0.0001596, -0.0001507, -0.0012035, -0.0268494, 0.1078350, 0.2952210, 0.3512440, 0.3037620, 0.1242870, 0.0076266, -0.0524563, -0.2097750, -0.4972090, -0.2121350, -0.0335701, -0.0404355, -0.1694020, -0.0712553, 0.0892602, -0.0703997, 0.0481584, 0.0232640, 0.0425058, 0.0682251, -0.0027273, -0.0760942, -0.0580954, -0.0011003, 0.0000712, -0.0027200, -0.0041817, -0.0319508, 0.0745275, 0.1690030, 0.1151090, 0.1101130, -0.1105660, 0.0214761, 0.0068199, -0.3813710, -0.2823210, -0.1673980, -0.1178200, -0.1324730, 0.1187530, 0.2890070, -0.0562912, -0.1198720, 0.0143165, -0.0609425, -0.0543038, 0.0103829, -0.0575157, -0.1382980, -0.0768722, -0.0127800, -0.0006663, -0.0013531, -0.0105394, -0.0456845, 0.0126631, 0.0457127, -0.1314480, -0.1630500, -0.0475870, -0.1486460, -0.2694510, -0.5406680, -0.2718570, -0.0732631, -0.0398482, 0.0100306, 0.2137620, -0.0334408, -0.0597591, -0.0259679, 0.2160890, 0.0246226, -0.0581974, -0.1031470, -0.1272830, -0.1592250, -0.1400030, -0.0246857, -0.0002617, -0.0002947, -0.0072413, -0.0737905, -0.1388600, -0.0205753, -0.1262140, -0.2031990, -0.0210511, -0.0872998, -0.3104650, -0.4189250, -0.0808216, 0.2419550, 0.2093200, 0.1344920, 0.2039580, 0.2056430, 0.0348242, 0.0875732, 0.2347530, 0.0496425, 0.0857716, -0.0954555, -0.0695400, -0.1075470, -0.0496879, -0.0060578, -0.0004823, 0.0000827, -0.0088316, -0.1073220, -0.1553890, -0.0603412, -0.0831358, -0.0903422, -0.0713940, -0.1012230, -0.3275170, -0.1007370, 0.2109270, 0.3590630, 0.2070610, 0.0029986, -0.0045322, 0.1302760, -0.0269694, 0.0385968, 0.1031730, 0.0285417, -0.0799988, -0.2015920, -0.1374340, -0.0655560, -0.0031629, -0.0043245, -0.0001153, 0.0001995, -0.0170580, -0.1335320, -0.1011350, -0.0134485, -0.0007464, -0.2739770, -0.3473840, -0.3029190, -0.2101100, 0.1070690, 0.4493450, 0.1838130, 0.1828000, 0.0121786, 0.0164507, 0.0658939, 0.0666135, -0.1030120, -0.0010587, 0.0509649, -0.1132840, -0.1944220, -0.0223606, -0.0486059, -0.0169642, -0.0000767, -0.0001917, 0.0005161, -0.0249294, -0.1530890, -0.1476500, -0.0637791, -0.0233529, -0.3859330, -0.2954080, -0.1061340, -0.0968597, 0.0469272, 0.1159590, 0.1768460, 0.2738600, 0.0959421, 0.0149073, 0.2013560, 0.1901570, -0.0212979, 0.0057110, -0.0310498, 0.0011483, -0.1456320, 0.0243401, 0.0058478, -0.0076824, -0.0004844, 0.0000655, -0.0004549, -0.0436790, -0.1322870, -0.1907830, -0.1192620, -0.1030090, -0.2479300, -0.2048930, -0.0193823, -0.0120534, 0.0850120, 0.0831677, 0.1112800, 0.1873970, 0.3026420, 0.2379210, 0.1311850, 0.0842144, -0.0474917, 0.0353648, -0.0458445, -0.0479299, -0.0403376, 0.0579451, 0.0278583, -0.0002652, -0.0003901, -0.0001813, 0.0004119, -0.0291408, -0.0350971, -0.1975410, -0.2500570, -0.1345970, -0.0443523, -0.0915601, 0.0494099, 0.0332545, 0.0308572, 0.2609820, 0.1667700, 0.1654720, 0.2080190, 0.0955515, 0.0300514, 0.0993713, -0.0822649, -0.0072415, -0.0561213, -0.0617550, 0.0063483, 0.0685819, 0.0524128, 0.0023324, -0.0003936, 0.0001821, 0.0004868, -0.0152645, -0.0297643, -0.1564980, -0.1541610, -0.0736406, -0.0901862, 0.1904020, 0.0382034, 0.0771217, 0.0835428, 0.0117179, -0.1339200, 0.1203610, 0.1289880, 0.0746762, 0.0143801, 0.0311340, 0.0636807, 0.0516620, 0.0067811, 0.0101712, 0.0843178, 0.0855225, 0.0219488, 0.0017015, 0.0001995, -0.0000835, 0.0003373, -0.0085061, -0.0282485, -0.0382453, -0.0016513, -0.0117173, 0.1580430, 0.1067470, 0.1527420, 0.0594140, 0.0057493, -0.0427738, 0.1382160, 0.1162080, 0.0995273, 0.0234769, 0.0950476, 0.1605760, 0.1163080, 0.0485142, 0.0599257, 0.0994014, 0.1219800, 0.0431443, -0.0016145, -0.0003230, 0.0002354, -0.0001093, -0.0000371, -0.0017496, 0.0010465, 0.0092050, 0.0170708, -0.0284947, 0.0330155, 0.0323313, 0.0098062, -0.1266870, -0.1269430, -0.1865320, -0.0623701, -0.0997912, -0.1067660, -0.0292704, 0.0714670, 0.1439590, 0.1340140, 0.0868582, 0.0996815, 0.0596227, 0.0407797, 0.0221418, -0.0001470, -0.0008585, 0.0005084, -0.0005770, 0.0000884, 0.0005450, 0.0003522, 0.0050672, 0.0237665, 0.0484253, 0.0564310, 0.0457916, 0.0392390, 0.0556246, 0.0783571, 0.0750730, 0.0090287, 0.0533879, 0.0408720, 0.0097442, -0.0256189, 0.0074334, 0.0456045, 0.0633217, 0.0583344, 0.0251658, 0.0027208, 0.0023866, 0.0000258, 0.0001390, -0.0002504, -0.0005616, 0.0003754, -0.0004834, -0.0001423, -0.0002497, -0.0007342, 0.0007615, 0.0111794, 0.0103772, 0.0011304, 0.0009501, 0.0034852, 0.0029721, 0.0005227, 0.0009948, -0.0029028, -0.0019260, -0.0014335, 0.0195874, 0.0222342, 0.0139028, 0.0009725, 0.0078494, -0.0022682, 0.0002367, 0.0000334, -0.0003047, 0.0004193, -0.0003548, -0.0002860, 0.0000064, 0.0002185, 0.0004969, -0.0003354, 0.0001833, 0.0001915, -0.0004099, 0.0001462, -0.0005908, 0.0000776, -0.0004455, 0.0001996, 0.0000880, 0.0001590, -0.0000095, 0.0000383, -0.0004437, 0.0001911, 0.0001864, -0.0001339, 0.0005391, 0.0000991, 0.0002011, -0.0002129, -0.0002318, -0.0001109, 0.0002367, -0.0003252, 0.0003481, -0.0004948, -0.0001932, 0.0001317, -0.0000433, 0.0002385, 0.0001812, -0.0002554, -0.0003207, -0.0015209, -0.0023757, -0.0012896, 0.0056042, -0.0042423, -0.0442124, -0.0195788, -0.0010814, -0.0007560, -0.0000044, 0.0007481, 0.0003333, -0.0000854, -0.0001021, 0.0009770, 0.0003437, 0.0001412, 0.0002652, 0.0006016, -0.0001461, -0.0001855, -0.0007798, -0.0002867, -0.0000725, -0.0005233, -0.0054681, -0.0120420, -0.0085665, -0.0104823, -0.0124457, -0.0235174, -0.0486661, -0.0450196, -0.0505519, -0.0303221, -0.0024257, -0.0122499, -0.0126460, -0.0101200, -0.0051022, -0.0046394, -0.0049501, -0.0019964, 0.0000857, 0.0000819, -0.0003183, -0.0004841, 0.0049260, 0.0011021, 0.0001265, -0.0012177, -0.0018132, -0.0017012, -0.0146968, -0.0341791, -0.0536658, -0.0497679, 0.0165960, -0.1525050, -0.2878260, -0.2120720, -0.2457950, -0.1802290, -0.1673100, -0.0824791, -0.0797042, -0.0393348, 0.0201118, -0.0736029, -0.0773892, 0.0467927, 0.0037407, 0.0001989, 0.0000635, -0.0000061, 0.0136154, 0.0026415, -0.0036421, -0.0121235, -0.0193062, -0.0437021, -0.0961928, -0.1738000, -0.1985950, -0.1047260, -0.0407430, -0.0406540, -0.1861520, -0.1549770, -0.1763300, -0.0670627, -0.0653862, -0.1711360, -0.1872460, -0.2293760, -0.1440760, -0.0059063, -0.0833067, 0.0253585, 0.0166754, -0.0042366, -0.0000293, 0.0001590, 0.0012060, -0.0011637, -0.0052096, -0.0144852, -0.0531817, -0.1142550, -0.2689250, -0.3132510, -0.2728860, -0.1261650, -0.0801579, -0.0797798, -0.1703120, -0.1940760, -0.2197700, -0.2150180, -0.2940480, -0.0688169, 0.0094561, -0.1546650, -0.0627190, -0.0513652, -0.0900252, -0.0467147, -0.0156481, -0.0061075, -0.0001837, -0.0004917, 0.0041999, -0.0007662, -0.0107624, -0.0408992, -0.0758604, -0.1758920, -0.3436330, -0.3505230, -0.2515790, -0.0626712, 0.0205728, -0.1080170, -0.1312610, -0.3128720, -0.2744630, -0.3104370, -0.1224060, -0.1474900, -0.1552890, -0.1299330, 0.0636646, 0.0953145, -0.0043587, 0.0041361, 0.0616519, 0.0041302, 0.0000128, -0.0034037, -0.0120268, -0.0070033, -0.0151183, -0.0323565, -0.0959255, -0.2143650, -0.3523460, -0.2453470, -0.1952190, -0.1138720, 0.0203138, 0.0869462, -0.0333729, -0.2594710, -0.0204865, -0.2626460, -0.1606830, -0.0220044, -0.0745273, 0.0461026, 0.1369850, 0.1695760, 0.0523245, 0.0061493, 0.0578545, 0.0002137, -0.0059831, -0.0020237, -0.0153059, -0.0124152, -0.0142673, -0.0193693, -0.0832555, -0.1878180, -0.2107440, -0.1963450, -0.2727040, -0.3110960, 0.0808106, 0.2324480, 0.1633320, -0.0205833, 0.0908851, 0.2064740, 0.1968160, 0.2063410, 0.1973320, 0.2157470, 0.1606340, 0.3332960, 0.3241340, 0.1014730, -0.0057400, 0.0009450, -0.0004468, -0.0013248, -0.0117890, -0.0193453, -0.0184266, -0.0852434, -0.1204750, -0.1786220, -0.1117860, -0.1470890, -0.1434990, -0.1100300, 0.0117189, 0.4479480, 0.4111080, 0.1772830, 0.1916600, 0.3708770, 0.4235210, 0.3564040, 0.0932284, 0.1988910, 0.2375410, 0.1115670, 0.1416600, 0.1555450, 0.0808490, 0.0068378, -0.0009098, 0.0000806, -0.0134264, -0.0293946, -0.0462819, -0.1400180, -0.1813020, -0.1176470, 0.1554230, 0.1525320, 0.1706920, 0.0054586, 0.0661914, 0.3357680, 0.2391590, 0.0117232, -0.1269620, -0.1080680, -0.0968496, 0.1111210, 0.1036120, 0.1551620, 0.0400101, 0.0252567, 0.1449960, 0.2716300, 0.0465459, 0.0004487, -0.0000301, -0.0033696, -0.0061519, -0.0237499, -0.0337262, -0.1570160, -0.2086170, -0.1459540, 0.0459151, 0.0311827, 0.0050628, -0.0173128, -0.0264561, 0.0334222, 0.1462330, -0.1248790, 0.0978735, -0.0865927, 0.0391026, 0.0382545, 0.1261790, 0.1261120, 0.0471239, 0.0955681, 0.1503940, 0.1390960, -0.0029518, -0.0009353, 0.0000236, -0.0009989, -0.0031347, -0.0194278, -0.0307216, -0.2086020, -0.1378410, 0.0673580, 0.1507850, 0.0821973, 0.0895311, 0.0922510, 0.0532563, 0.2411150, 0.2873330, 0.1762980, 0.1905050, 0.0750578, -0.1139850, -0.1601860, -0.0306676, -0.1503280, -0.2527370, -0.1267160, -0.0794325, 0.0362791, 0.0150438, -0.0021140, 0.0001794, -0.0001658, -0.0058738, -0.0145068, -0.0397892, -0.0903721, -0.0297901, 0.0862981, 0.0165181, 0.1833150, 0.1003500, 0.0535214, 0.1559950, 0.1385990, 0.3186370, 0.1471820, 0.1135970, 0.0513413, -0.3194850, -0.2999160, -0.2599480, -0.2768500, -0.3751920, -0.2768700, -0.0869781, 0.0046037, -0.0115697, -0.0017453, 0.0011291, -0.0001582, -0.0006243, -0.0082537, -0.0105418, -0.0103123, -0.0737406, -0.0860318, -0.0448330, 0.0628199, 0.0985789, -0.0949665, -0.0755376, 0.0064643, 0.1917320, 0.1076300, -0.0055020, -0.1710480, -0.2170950, -0.2383860, -0.2630510, -0.2796330, -0.2614400, -0.1769220, -0.0277394, -0.0171374, -0.0073907, -0.0003372, 0.0003913, 0.0000389, 0.0005934, -0.0013943, -0.0091408, -0.0141913, 0.0122404, -0.0174038, -0.0140048, 0.0558147, 0.1233700, 0.0204230, 0.1446730, 0.0872187, 0.2241730, -0.0908745, -0.1010340, -0.2420740, -0.1619290, -0.2318780, -0.3218430, -0.3361010, -0.2789330, -0.1304060, -0.0649746, 0.0064592, -0.0068021, -0.0043617, -0.0002806, -0.0004941, -0.0024479, -0.0136082, -0.0716647, 0.0404136, 0.0069666, -0.0845680, 0.0260834, -0.0929246, 0.0199991, 0.1286390, 0.1031420, 0.1957420, 0.1721380, -0.2871130, -0.2631310, -0.2509340, -0.1209920, -0.1578000, -0.2742370, -0.2321120, -0.2043440, -0.1727040, -0.0387348, 0.0078355, -0.0165159, -0.0051042, 0.0004650, -0.0002990, -0.0045724, -0.0468792, -0.1032550, -0.0297552, 0.0208269, -0.0963395, -0.1409190, 0.0323368, 0.1469670, 0.2099680, 0.0266931, 0.1964550, 0.2201820, -0.1993870, -0.2432850, -0.2511510, -0.1534650, -0.2339740, -0.2068970, -0.2694310, -0.1654660, -0.1147730, -0.0412602, 0.0125038, -0.0086431, -0.0050007, -0.0011171, -0.0000708, -0.0027699, -0.0885954, -0.1522080, -0.1635250, -0.0949685, 0.0241995, -0.0847913, -0.0263771, -0.1625810, 0.1301600, 0.0551596, 0.1698680, 0.2374230, -0.3473520, -0.4896300, -0.1972570, -0.1688950, -0.2012030, -0.1078770, -0.2609420, -0.1857590, -0.1052240, -0.0308230, 0.0421046, 0.0052817, 0.0046801, 0.0008176, -0.0002676, -0.0031039, -0.1114500, -0.1316460, -0.1450860, -0.0556837, 0.0405407, 0.0406133, -0.1468610, -0.2209740, -0.2990960, -0.1132320, 0.2289940, -0.0226767, -0.1651470, -0.2031210, -0.2351130, -0.1728370, -0.0826143, -0.2671690, -0.3202650, -0.1625250, -0.0648593, 0.0188142, 0.0520590, 0.0026561, 0.0032873, 0.0003423, 0.0002525, -0.0093615, -0.1490130, -0.1697400, -0.1275940, 0.0617709, -0.0131870, 0.0327358, -0.1229370, -0.2669360, -0.1524040, -0.0341451, -0.0155686, 0.1107770, 0.0362067, -0.0022122, -0.0599504, -0.1007240, -0.0458326, -0.1671910, -0.2483460, -0.1237740, -0.0484088, 0.0262832, 0.0333477, 0.0035459, -0.0004568, 0.0000831, -0.0001509, -0.0082042, -0.1311310, -0.1576990, -0.1614790, -0.0983464, -0.0271603, -0.2146130, -0.1204780, -0.0511185, -0.0102367, -0.0172797, -0.0086106, 0.0356862, -0.0008109, -0.1037240, -0.1387040, -0.0042489, -0.0450212, 0.0549939, -0.1052110, -0.1171830, -0.0338309, 0.0370854, 0.0084509, -0.0005685, 0.0004985, 0.0001391, 0.0004042, -0.0066971, -0.0208325, -0.0541832, -0.0545460, -0.0279622, 0.0861729, -0.0238228, 0.0701247, 0.0688581, 0.0677333, -0.0003010, -0.0273165, -0.0712901, -0.2043550, -0.0447297, 0.1108890, 0.0701997, -0.0574947, 0.0398716, -0.0752669, -0.0867406, 0.0010814, 0.0105654, 0.0005186, 0.0019751, 0.0004898, 0.0000783, 0.0000880, -0.0051666, -0.0029098, -0.0163025, 0.0371789, 0.0462296, 0.1819420, 0.1725390, 0.2437020, 0.2466810, 0.1341670, 0.2134740, 0.0204412, -0.0435006, -0.0741459, 0.0482166, 0.1687530, -0.0374622, -0.0825204, -0.0194244, -0.0908508, -0.0510673, -0.0006060, 0.0138643, 0.0045058, 0.0019314, 0.0000433, -0.0000366, 0.0005653, -0.0014824, -0.0081934, -0.0288359, -0.0450214, -0.1340890, 0.0043790, 0.0818007, 0.1067300, 0.1088680, -0.0423901, -0.0698845, -0.0731049, -0.1756890, -0.0842703, -0.2311330, -0.0108722, -0.0339751, -0.0192098, -0.0497039, -0.0527932, -0.0218753, 0.0255501, 0.0131684, -0.0021646, -0.0014473, 0.0003837, 0.0003329, -0.0002340, -0.0001996, 0.0000147, -0.0214468, -0.0440393, -0.1035470, -0.0814558, -0.0826587, -0.1012190, -0.1470570, -0.1260050, -0.1349200, -0.0332325, -0.0786821, -0.0501752, 0.0115944, -0.0093840, -0.0259576, -0.0216663, 0.0099186, 0.0088069, 0.0114468, 0.0222694, 0.0111649, -0.0012783, -0.0011246, -0.0004241, 0.0005031, -0.0002972, -0.0005202, -0.0000920, -0.0032916, -0.0110813, -0.0164502, -0.0214685, -0.0195509, -0.0274302, -0.0232062, 0.0089620, 0.0127414, -0.0136233, 0.0126728, 0.0560671, 0.0218311, -0.0492376, -0.0583642, 0.0106858, 0.0098422, -0.0028383, -0.0032529, 0.0000203, -0.0001610, 0.0002747, -0.0003642, 0.0000233, 0.0003888, -0.0004667, -0.0002064, -0.0006537, -0.0000169, -0.0002388, 0.0013627, 0.0048464, 0.0029864, -0.0011811, -0.0027849, -0.0057855, -0.0064123, -0.0202523, -0.0044386, 0.0094814, -0.0008311, -0.0083774, -0.0010512, 0.0009307, 0.0011105, -0.0062498, -0.0035503, 0.0000050, 0.0006124, 0.0001834, 0.0007352, -0.0003356, 0.0001669, 0.0002735, 0.0005575, 0.0005520, -0.0003746, 0.0001114, 0.0002434, -0.0002089, -0.0005329, -0.0002569, 0.0001482, 0.0007505, -0.0009711, -0.0016757, -0.0009428, 0.0000090, -0.0000003, 0.0001438, -0.0000234, 0.0000752, 0.0003098, 0.0001745, -0.0003846, 0.0000537, -0.0004893, -0.0002440, 0.0001797, -0.0005552, 0.0000238, -0.0002685, -0.0000674, 0.0003284, -0.0002478, 0.0001471, -0.0029606, -0.0047485, -0.0039611, -0.0013322, -0.0061919, -0.0114533, -0.0163846, -0.0196935, 0.0288580, 0.0079651, -0.0217685, -0.0197838, -0.0184318, -0.0234417, -0.0161470, -0.0043655, -0.0052166, -0.0053010, -0.0003120, -0.0003158, -0.0004724, -0.0000321, -0.0001589, -0.0004007, -0.0005902, -0.0011178, -0.0006807, 0.0000975, -0.0052272, -0.0177895, -0.0301389, -0.0530679, -0.0679688, -0.0928143, -0.0671340, -0.0201530, -0.1160630, -0.0928708, -0.0982139, -0.0922614, -0.0915556, -0.0581269, -0.0870196, -0.0829766, -0.0364480, -0.0449873, -0.0240138, -0.0046095, 0.0005302, 0.0002785, 0.0002095, -0.0001340, 0.0063203, -0.0025565, -0.0046587, -0.0213588, -0.0870220, -0.0500159, -0.1388840, -0.2730460, -0.0577059, -0.0919013, -0.0963682, -0.1817150, -0.1490310, -0.0635236, -0.0728023, 0.0568308, 0.0374945, -0.0868734, -0.0075471, -0.1323670, -0.0760290, -0.0784149, -0.0439079, -0.0015082, -0.0056411, 0.0000889, 0.0000352, 0.0001284, 0.0214753, 0.0079800, -0.0317171, -0.0508681, -0.0849246, -0.0871480, -0.2046240, -0.2373780, -0.1729080, 0.0020284, 0.0105580, 0.0529734, 0.1102410, 0.2237850, 0.0390340, -0.0656993, 0.0042876, -0.0869904, 0.0779894, 0.1887010, 0.1218390, 0.0890131, 0.1108760, 0.0121808, -0.0042155, -0.0032545, -0.0000518, 0.0000442, -0.0002819, 0.0142249, -0.0660512, 0.0670777, 0.0021106, -0.0368286, -0.1266830, -0.1188450, -0.0212096, 0.1414860, 0.0374128, 0.0256343, 0.0875506, 0.1728610, 0.0366399, 0.0787355, 0.0786726, 0.0742944, 0.0660241, 0.1693900, 0.1858790, 0.0556740, 0.0701350, 0.0105959, -0.0081418, -0.0045246, -0.0002752, -0.0002502, 0.0036072, -0.0072517, -0.0604412, 0.0860831, 0.0610521, 0.0828237, 0.1078860, 0.0526612, 0.1912060, 0.0398774, 0.0718703, -0.0391114, 0.1780010, 0.1441340, 0.2217390, 0.2346040, 0.2907970, 0.3101140, 0.5119680, 0.3392910, 0.2836920, 0.2477690, 0.0568807, -0.0465601, 0.0224611, -0.0007248, -0.0000225, 0.0000780, 0.0006528, 0.0412993, -0.0289122, 0.1924010, 0.2022800, 0.1502550, 0.0047822, 0.0521477, 0.0283685, -0.0453293, 0.2174480, 0.2077000, 0.2729680, 0.0834219, 0.3267660, 0.2566410, 0.3595640, 0.4912040, 0.4017180, 0.3339780, 0.4860400, 0.4670430, 0.0492704, -0.0937535, 0.0738914, -0.0011544, -0.0002733, 0.0000343, 0.0045402, 0.0440144, -0.0063680, 0.1624760, 0.1768090, 0.0276400, -0.0708388, -0.0862770, -0.1937800, 0.0186575, 0.2022280, 0.0156261, 0.0186780, 0.1705750, 0.0300026, 0.1249650, 0.3554900, 0.1249990, 0.0112048, 0.1637330, 0.3368660, 0.3214750, 0.2084440, 0.1104160, 0.0243618, -0.0064017, 0.0000769, 0.0031102, 0.0052412, 0.0198471, -0.0037514, 0.1060140, 0.1529820, -0.0001329, -0.0188449, -0.0529183, 0.0871545, 0.1444580, 0.0724872, 0.0394897, -0.1533680, 0.0539265, -0.0532534, 0.0268513, 0.0525686, 0.0238707, -0.0797106, 0.1329200, 0.1044740, 0.2416860, 0.1122930, 0.1712070, 0.0698287, 0.0476753, -0.0004504, 0.0000574, 0.0249519, 0.0453466, -0.0260457, 0.0073399, -0.0729200, -0.0702917, -0.0271144, 0.0822278, 0.2034580, 0.1561600, 0.2199980, 0.1730230, 0.0589749, 0.1351760, 0.1262310, 0.0213891, 0.1042320, 0.2001770, 0.0410100, 0.0626250, 0.2295290, 0.1609270, 0.0944629, 0.2322300, 0.0425292, 0.0151979, 0.0002034, 0.0004280, 0.0361657, 0.0345683, 0.0226698, 0.0044187, -0.0717448, -0.0329337, 0.0768524, 0.0193971, 0.3226390, 0.1406180, 0.1561700, 0.1304910, 0.1012710, 0.3179370, 0.0962799, 0.1510970, 0.0622099, 0.0440708, -0.0385291, 0.0506512, 0.0489516, 0.0045396, -0.0260964, 0.0175931, 0.0371339, 0.0051066, -0.0000893, 0.0009856, 0.0329986, 0.0346019, 0.0286120, -0.0639779, -0.0307336, 0.0305482, 0.1168930, 0.1526180, 0.1701940, -0.0494586, 0.0592643, 0.1397220, -0.0117081, 0.2309080, -0.0661800, 0.0453053, 0.0609023, -0.0448203, 0.0295151, -0.0534656, -0.0653482, -0.1193590, -0.1045000, -0.0068110, 0.0587157, 0.0102376, 0.0003796, 0.0017325, 0.0045293, -0.0150024, 0.0369559, -0.0983804, 0.0062510, 0.0950384, 0.1154240, 0.1335670, 0.0176851, -0.0482909, -0.1033890, -0.3015750, -0.0731507, 0.0551170, -0.2355630, 0.1696420, -0.0863696, -0.1581480, 0.0435400, -0.1300370, -0.0820036, -0.3796090, -0.2007100, -0.0197187, -0.0259482, -0.0165629, 0.0000103, 0.0008169, 0.0016594, -0.0554908, 0.0255480, 0.0227034, -0.0234169, -0.0111197, -0.0624799, -0.1861210, -0.2399330, -0.1249530, -0.0671551, -0.2726620, -0.0823410, -0.0649191, -0.0890281, 0.3565870, -0.1517150, 0.0336144, -0.0451081, -0.2187230, -0.2959850, -0.1513930, -0.0735502, -0.1003100, -0.0600352, -0.0016583, -0.0002955, 0.0005966, -0.0209624, -0.0903838, 0.0315293, 0.0407880, -0.0537760, 0.0474117, 0.0660972, 0.0617333, 0.0588900, -0.0326165, 0.0446945, -0.3871070, -0.2170090, -0.0549052, 0.0302025, 0.2141970, -0.0512684, -0.1957730, -0.2060420, -0.1325320, -0.0337154, 0.0739022, -0.0870623, -0.1183230, 0.0095515, -0.0152735, 0.0002921, 0.0005765, -0.0489984, -0.0714102, -0.0027376, -0.0482412, -0.2401710, -0.0065051, 0.1801930, 0.0241316, 0.0168819, -0.1868140, 0.0634771, -0.0701605, -0.3624710, -0.0784074, -0.0142766, -0.2044080, -0.2195220, -0.2011210, -0.1026430, -0.1749950, -0.1110630, 0.0321907, -0.1229520, -0.1941180, -0.0956950, -0.0239755, 0.0005241, -0.0001971, -0.0570210, -0.0608282, 0.0269282, 0.0813918, -0.0851498, -0.0298262, -0.0972515, 0.0737680, -0.1664160, -0.2313200, -0.0392215, -0.0112815, 0.0937930, 0.0421086, -0.1674180, -0.3172890, -0.1879600, -0.0925224, -0.1627870, -0.1467790, 0.0784447, 0.1996690, -0.0223590, -0.1625450, -0.0028755, -0.0110289, -0.0002032, -0.0003655, -0.0102785, -0.0238524, 0.0142510, 0.0543664, 0.0162166, -0.1915260, 0.0141058, 0.1459560, -0.1329260, 0.0756334, -0.1844400, 0.0005771, 0.0272074, -0.0483295, -0.2196240, -0.3403230, -0.1274690, -0.1320410, 0.0228081, -0.0194635, -0.0148039, -0.1398030, -0.1572530, -0.1471420, 0.0174312, -0.0083748, 0.0000543, 0.0026997, 0.0079020, 0.0585969, 0.0596139, 0.0207107, -0.0651435, -0.0698725, 0.0687001, 0.0991084, -0.1353530, -0.2239450, -0.1412200, 0.0758037, -0.2040840, -0.2828420, -0.1508180, -0.1572590, -0.0308807, 0.0008230, -0.1076440, -0.0482908, -0.1916730, -0.3124110, -0.1352300, -0.0742711, -0.0177354, -0.0004364, -0.0004856, 0.0051093, 0.0044783, 0.0254083, 0.0988495, 0.0293241, 0.1476330, -0.1145290, 0.0161749, -0.0053503, -0.3159660, -0.2583660, -0.1851950, -0.0599630, -0.1949490, -0.2199790, 0.0633933, 0.0761139, -0.1330090, 0.1766430, 0.0267224, 0.0075890, -0.0654009, -0.0780130, -0.1259500, -0.0326499, -0.0098455, 0.0001412, -0.0001793, -0.0004608, -0.0057715, -0.0015625, 0.0529051, 0.2001410, 0.0433474, -0.1217850, -0.0831392, 0.0210711, -0.2088990, -0.1304140, -0.1752290, -0.3164390, -0.1900840, 0.0606879, 0.0593017, 0.0532902, 0.0567409, 0.2510280, 0.2920820, 0.2733790, 0.1161130, 0.0110458, 0.0288635, 0.0344372, 0.0000953, -0.0002243, -0.0002278, -0.0000593, -0.0028079, -0.0076194, 0.0680342, 0.0889109, 0.1139380, 0.1208830, 0.1831630, 0.0054352, -0.0645382, 0.2087710, 0.2558040, 0.1876470, 0.4296460, 0.2404240, 0.2757220, 0.3780520, 0.3619630, 0.4232380, 0.2838970, 0.2795690, 0.1421610, 0.1037170, 0.0826038, 0.0676764, 0.0164258, 0.0001049, 0.0001738, -0.0001649, -0.0004613, 0.0011719, 0.0610449, 0.0782030, 0.1258700, 0.2248690, 0.3088080, 0.4007980, 0.3899200, 0.4059530, 0.5247850, 0.5900680, 0.5998030, 0.6303070, 0.5858590, 0.5318920, 0.3259150, 0.1818500, 0.1136030, 0.0901249, 0.0381817, 0.0996187, 0.0700663, 0.0585422, 0.0093310, 0.0004610, 0.0000549, 0.0000874, 0.0042533, 0.0138563, 0.0368507, 0.0885163, 0.1091620, 0.1373660, 0.1569530, 0.3141470, 0.2217040, 0.3011910, 0.3517700, 0.3948850, 0.3547420, 0.3170630, 0.2132630, 0.1711600, 0.0627690, 0.0639051, 0.0974874, 0.0736183, 0.0187953, 0.0045967, -0.0187689, -0.0033602, -0.0010070, -0.0005062, 0.0000042, 0.0003116, -0.0002392, 0.0026591, 0.0050781, 0.0193732, 0.0185389, 0.0368493, 0.0686480, 0.1014510, 0.0146300, 0.0394384, 0.0394747, 0.1125430, 0.0675983, 0.1270280, 0.0965207, 0.0061421, -0.0093343, 0.0219235, 0.0435220, -0.0055314, -0.0122110, -0.0071703, -0.0104459, -0.0006509, -0.0002580, 0.0002702, -0.0001126, -0.0000569, -0.0006562, 0.0001234, 0.0000212, -0.0012942, 0.0017243, 0.0072002, 0.0164888, 0.0227988, 0.0164188, 0.0055359, -0.0003847, 0.0074301, -0.0081029, 0.0078767, 0.0013703, -0.0185771, -0.0425132, -0.0449022, -0.0271393, -0.0191053, -0.0050290, -0.0036768, -0.0005833, 0.0000710, -0.0000958, 0.0002850, 0.0002602, -0.0003957, 0.0002776, -0.0005238, 0.0003161, 0.0002342, -0.0010499, -0.0047776, -0.0045362, 0.0011804, 0.0051668, 0.0008035, -0.0023329, 0.0010897, -0.0067325, 0.0001788, 0.0001458, -0.0002862, -0.0073150, -0.0060303, -0.0006131, 0.0035916, -0.0019791, 0.0015724, -0.0000859, -0.0002300, 0.0001845, 0.0002142, 0.0001693, 0.0002562, -0.0004886, 0.0002208, -0.0000615, -0.0002446, 0.0006200, -0.0006892, 0.0003035, 0.0001429, 0.0002405, -0.0001706, -0.0000409, 0.0008100, -0.0002894, 0.0002721, 0.0000997, 0.0000932, 0.0000652, -0.0003129, 0.0000574, -0.0003328, -0.0005217, -0.0000424, 0.0000119, 0.0002876, -0.0000030, -0.0002891, 0.0002511, -0.0003220, -0.0001238, 0.0006660, 0.0000305, 0.0004333, 0.0057587, 0.0086845, 0.0050045, 0.0020963, 0.0059541, 0.0041029, 0.0030876, 0.0045901, -0.0083433, 0.0066455, 0.0089444, 0.0073616, 0.0051845, 0.0041125, 0.0027377, 0.0016763, 0.0005983, 0.0002596, -0.0001970, 0.0000016, -0.0000049, 0.0004436, -0.0001712, 0.0000738, 0.0002726, -0.0004850, 0.0001729, 0.0004534, 0.0032130, 0.0137701, 0.0230537, 0.0137429, 0.0162196, 0.0331596, 0.0197100, -0.0465653, -0.0320950, 0.0234085, 0.0619786, 0.0501229, 0.0382313, 0.0184501, 0.0100447, -0.0074126, -0.0072689, 0.0023674, -0.0006861, -0.0008047, 0.0000696, 0.0004588, -0.0005403, 0.0000609, 0.0002182, -0.0001757, 0.0046954, 0.0385774, 0.0531435, 0.0705921, 0.0561886, 0.0412068, -0.0072541, -0.0190750, 0.0203342, -0.0925318, -0.0675388, 0.0380230, 0.0143048, 0.0501671, 0.1104770, 0.1018750, 0.0641680, 0.0242579, 0.0258098, 0.0399808, 0.0209005, -0.0000514, 0.0009222, 0.0006360, -0.0002151, 0.0002420, -0.0004620, -0.0001262, 0.0050639, 0.0429948, 0.0123631, 0.0197022, 0.0675787, -0.0287385, 0.0608246, -0.0254154, 0.0063061, -0.0064079, 0.0629591, 0.1711170, 0.1712290, 0.0204857, 0.0390461, 0.1148140, 0.0591404, 0.1266720, -0.0016371, 0.0004337, 0.0097077, -0.0023792, -0.0001976, 0.0002380, 0.0000254, -0.0006167, 0.0002963, -0.0036581, -0.0093664, 0.0083689, -0.0042169, 0.1464060, 0.1085410, 0.0524516, 0.0511712, -0.0389431, 0.0052386, -0.1793310, -0.0270406, -0.0484835, 0.0198680, 0.0153419, 0.0237381, 0.1114840, 0.1499830, 0.1386460, 0.0840131, 0.0838488, 0.0230840, 0.0097781, 0.0039590, 0.0019812, 0.0000734, 0.0001388, -0.0018165, -0.0151561, -0.0060773, -0.0205855, 0.0028295, 0.0893538, 0.0946388, 0.1634670, 0.0514631, 0.0393133, 0.1849240, 0.0420416, 0.0529174, 0.0354609, 0.0220129, 0.0849720, 0.0787137, 0.0192670, -0.0331179, 0.0195109, -0.0231885, -0.0157252, 0.0498236, 0.0446821, 0.0165288, 0.0066221, 0.0001192, 0.0012189, -0.0059696, -0.0201363, -0.0382119, -0.0122622, -0.0885509, 0.0015494, 0.1416350, 0.0874939, 0.0134702, -0.1141290, -0.1692130, -0.1365860, 0.1340720, 0.0915576, 0.1928550, 0.1185490, 0.0201770, -0.0481314, -0.0365590, -0.0998683, -0.0426324, -0.0918874, -0.0083167, -0.0027568, 0.0139270, 0.0013728, -0.0007355, 0.0004967, -0.0265288, -0.0331346, -0.0630802, -0.0100658, -0.0379844, 0.1261310, 0.0587783, 0.0721450, 0.0382138, 0.0980791, 0.0349031, 0.1323140, 0.0098041, 0.1660560, -0.0256453, -0.0181765, -0.0991081, 0.0696598, 0.0246993, -0.0947410, 0.0328029, -0.0032167, 0.0284309, 0.0556794, 0.0019981, 0.0008053, 0.0002685, 0.0002248, -0.0186900, -0.0461767, -0.0997624, -0.0692614, 0.0666496, 0.1677080, 0.0726704, 0.0111229, -0.0087746, 0.1434480, 0.2090280, 0.0115815, 0.1429870, 0.1685720, 0.1964370, -0.0313534, -0.1355280, -0.1919540, -0.2207690, -0.0937354, 0.0919762, -0.0857582, 0.0044370, 0.0660708, 0.0106482, 0.0001005, -0.0003517, -0.0019092, -0.0245337, -0.0409008, -0.1178210, -0.0855774, 0.0637723, -0.0895092, 0.0216964, 0.0824533, 0.1261150, -0.0620473, 0.0549855, 0.2165920, 0.2227560, 0.2376930, 0.2139940, -0.0316107, -0.2474920, -0.1172210, -0.0810773, -0.1817840, -0.3676800, -0.2165710, 0.0371294, 0.0563601, 0.0262172, 0.0003845, 0.0000850, -0.0034487, -0.0103019, -0.0138975, -0.0566165, -0.0158256, -0.0728674, -0.2025300, -0.0568224, 0.0195501, 0.0441236, 0.0777037, 0.0650075, 0.0709896, 0.2738570, 0.4584440, 0.5809590, 0.1828880, -0.1462170, -0.1422880, -0.2364430, -0.1862540, -0.2598380, -0.1715230, 0.0260478, 0.0486485, 0.0329940, 0.0012029, 0.0000710, -0.0021913, -0.0030886, -0.0178669, -0.0963547, -0.1111310, -0.1691930, -0.0353621, 0.0174058, 0.0842942, 0.0608142, 0.0732645, -0.0944976, -0.0801339, 0.2374620, 0.6025200, 0.7300970, 0.3165530, -0.0367017, -0.2067120, -0.0947194, -0.1851860, -0.2185560, -0.2191460, -0.1012520, 0.0187088, 0.0208933, 0.0002485, 0.0000311, -0.0004197, 0.0012681, 0.0243599, -0.1705730, -0.1591610, -0.2119860, -0.1850260, -0.0897955, -0.0162946, -0.0328595, -0.0569722, -0.1150210, 0.0236759, 0.1828050, 0.5753930, 0.8545570, 0.1512090, -0.2102400, -0.2422400, -0.0351212, -0.2723380, -0.2391410, -0.1359280, -0.0800782, -0.0406415, 0.0019721, -0.0022514, -0.0000059, 0.0015819, 0.0023730, 0.0402589, -0.0015318, -0.1413910, -0.1635200, -0.2233960, -0.1552460, -0.0124880, -0.0463415, -0.1138710, -0.1834580, -0.0279555, 0.1001860, 0.5491420, 0.7741890, 0.1805190, -0.3923550, -0.2794340, -0.1997950, -0.1594340, -0.1389060, -0.0783957, -0.0981680, -0.0444254, -0.0201681, 0.0001152, 0.0005006, 0.0028056, 0.0075902, 0.0490354, 0.1880040, -0.0426678, -0.0452289, -0.1012180, -0.0526180, -0.1268610, -0.1778440, -0.1885840, -0.2080960, 0.0697381, 0.2495580, 0.6787270, 0.6746890, 0.0197272, -0.4537340, -0.3454470, -0.1453210, -0.0923663, -0.1516940, 0.0302579, -0.0516196, -0.0233983, -0.0412566, -0.0024563, -0.0002781, 0.0014707, 0.0171171, 0.1093190, 0.0790923, 0.0142729, -0.0455121, -0.0558546, 0.0159821, 0.0811971, -0.0601906, -0.2309610, -0.0625144, 0.2929020, 0.5692500, 0.6251120, 0.2969540, -0.4111060, -0.4905320, -0.1424500, -0.2067100, -0.1816030, -0.0367363, 0.1633560, 0.0037986, -0.0098893, -0.0296042, -0.0064593, -0.0004703, 0.0002948, 0.0207687, 0.1259970, 0.0403144, 0.0532138, -0.0545104, -0.0366236, -0.0178235, -0.0088144, -0.0439925, -0.0659713, 0.1266210, 0.3173910, 0.4602050, 0.3429760, -0.1258380, -0.4839980, -0.2835080, -0.0731216, -0.0347764, -0.0899840, -0.0197937, 0.1568790, -0.0410240, -0.0649900, -0.0168807, -0.0168695, -0.0002863, -0.0001562, 0.0172252, 0.1580280, 0.0782566, 0.0783170, -0.0750648, -0.0737261, -0.0536284, -0.1180700, -0.0602432, 0.0172440, 0.4033200, 0.4047380, 0.3195440, 0.0460024, -0.3054360, -0.3290080, -0.2521520, -0.0836554, -0.0797597, 0.0316627, -0.0620076, 0.0347180, -0.0383244, -0.0071945, -0.0028442, -0.0009598, 0.0002928, -0.0006067, 0.0187688, 0.1365470, 0.1083550, -0.0092669, -0.0977838, -0.1914070, -0.1179190, -0.0080103, 0.0393971, 0.1175210, 0.2253860, 0.2426770, -0.0133679, -0.1956190, -0.1442300, -0.0592671, -0.1682280, -0.1547690, 0.0162351, -0.0609491, -0.0719075, -0.0023166, -0.0065952, 0.0170917, -0.0053192, -0.0007390, 0.0002669, -0.0020631, 0.0043043, 0.0239064, 0.0549161, -0.2290350, -0.0875590, -0.0002974, 0.0221951, 0.1025840, 0.1294620, 0.1116410, 0.0554162, 0.0052760, 0.0772327, 0.0311995, -0.1113770, -0.0488043, -0.0298491, -0.2508240, -0.0080795, -0.1065890, -0.0048443, -0.0096286, -0.0613693, 0.0002711, -0.0019091, 0.0003867, -0.0000925, 0.0004213, -0.0203694, -0.0555881, 0.0480952, -0.1537080, -0.1776640, 0.0368231, 0.1085020, 0.2169580, 0.0992585, 0.0148041, -0.1345630, -0.0252074, 0.0352268, -0.0709905, -0.1873790, -0.0315203, 0.0169304, -0.1178940, 0.0276422, 0.0069333, -0.0722941, -0.0813994, -0.0955522, 0.0118173, -0.0012700, -0.0002159, -0.0000314, 0.0004618, -0.0099167, -0.0027493, 0.0558792, -0.0157474, -0.1161880, 0.0122477, 0.0513413, -0.0503886, 0.0522681, 0.0477631, -0.0224891, 0.1221950, 0.0456912, -0.0512559, -0.0529112, -0.0921731, -0.0223287, 0.0324134, 0.0164797, -0.0162554, -0.0867037, -0.0910200, -0.0844393, -0.0212856, 0.0022995, 0.0000632, 0.0003542, 0.0000602, 0.0038479, 0.0348487, 0.0970150, 0.0697997, -0.0389306, -0.0223672, -0.0401229, 0.0644562, 0.0040990, -0.0640102, -0.0106529, 0.1293660, -0.1463890, -0.1149340, -0.0066140, -0.0669290, -0.0194815, 0.0576524, 0.0403378, 0.0282854, -0.0280634, -0.0400779, -0.0357252, 0.0025995, 0.0023443, 0.0001769, 0.0002737, -0.0000737, 0.0012159, 0.0068535, 0.0289482, 0.0433478, 0.0344849, 0.0631877, -0.0785552, -0.2295210, -0.0602180, 0.0177678, 0.0137277, 0.0743199, -0.0459431, -0.0824584, 0.0301426, 0.0054933, 0.0120562, 0.0449685, -0.0385825, -0.0131766, -0.0045548, 0.0024849, 0.0155616, -0.0031606, 0.0001296, 0.0001488, 0.0001505, -0.0002110, 0.0003758, -0.0005037, 0.0034859, 0.0030785, -0.0060265, 0.0394902, 0.0261420, -0.0129471, 0.0793803, 0.0672223, 0.1027640, 0.1469460, -0.0324774, 0.0001034, 0.0355904, 0.0441849, -0.0196888, 0.0214635, 0.0161073, -0.0135914, 0.0213774, 0.0312630, 0.0213697, -0.0008556, 0.0002008, 0.0005436, 0.0000020, 0.0000089, 0.0000546, -0.0002612, 0.0001789, -0.0171876, -0.0277109, -0.0399350, -0.0363105, -0.0408693, 0.0071178, 0.0405383, -0.0210690, 0.0039320, -0.0096018, 0.0355123, -0.0023356, -0.0386908, -0.0343865, 0.0127348, -0.0142573, -0.0469396, -0.0148005, -0.0003149, -0.0013905, -0.0004852, -0.0001175, -0.0002495, 0.0001352, 0.0004917, -0.0003260, -0.0002153, 0.0000667, -0.0000035, 0.0003664, -0.0051303, -0.0055264, -0.0017198, -0.0010384, -0.0042851, -0.0045996, -0.0161431, -0.0220508, -0.0156749, -0.0151816, -0.0203522, -0.0382230, -0.0140321, -0.0074339, -0.0120837, -0.0046893, 0.0009547, 0.0000281, 0.0001688, 0.0001548, -0.0005054, -0.0000853, -0.0002870, 0.0005977, -0.0002801, -0.0008289, 0.0002485, -0.0002610, -0.0001925, 0.0001459, -0.0000918, 0.0002065, -0.0000703, -0.0016892, -0.0009004, 0.0001026, -0.0000871, 0.0000966, -0.0001143, 0.0000033, -0.0006902, -0.0002631, -0.0002573, 0.0001620, 0.0000060, -0.0005478, -0.0000222, -0.0001621, -0.0000668, 0.0000886, 0.0001062, -0.0002104, -0.0002561, 0.0003549, 0.0000893, -0.0004135, -0.0004071, 0.0007590, 0.0015954, 0.0023245, 0.0052207, 0.0075119, 0.0086987, 0.0007425, 0.0157851, 0.0533222, 0.0240942, -0.0026639, -0.0016622, -0.0019426, -0.0049756, -0.0011286, -0.0002642, -0.0000905, 0.0001473, 0.0001179, 0.0001904, 0.0003844, 0.0000271, 0.0000608, 0.0001996, 0.0006455, -0.0003671, -0.0013115, -0.0028631, -0.0054180, -0.0082921, 0.0031770, 0.0014916, -0.0056295, -0.0582773, -0.1055550, -0.1101050, -0.0625213, -0.0663812, -0.0526480, -0.0501678, -0.0444139, -0.0361615, -0.0208184, -0.0080685, 0.0005489, 0.0026550, -0.0002504, -0.0000648, -0.0003980, 0.0003987, -0.0000277, -0.0000142, -0.0006268, -0.0172481, -0.0263826, -0.0386434, -0.0252749, -0.0107826, -0.0097460, 0.0287034, 0.0449523, -0.0293881, -0.0923367, -0.1566450, -0.0940894, -0.0956575, -0.2156630, -0.2303630, -0.1457640, -0.0834702, -0.0560080, -0.0533479, -0.0236226, 0.0121857, 0.0021270, -0.0001774, 0.0002620, -0.0001519, 0.0006852, 0.0003905, -0.0053403, -0.0321107, -0.0171726, -0.0254270, -0.0415727, -0.0331705, -0.1074290, 0.0119977, -0.0744164, -0.1718120, -0.1649640, -0.0712685, -0.2643310, -0.0966607, -0.1123720, -0.2120310, -0.1275890, -0.1121110, -0.0466199, -0.0513849, -0.0502339, -0.0022138, 0.0067795, -0.0011619, 0.0002975, 0.0001891, 0.0000232, 0.0006851, -0.0069324, -0.0156352, -0.0167919, -0.0215715, 0.0361687, -0.0419178, -0.0973307, 0.0786042, -0.0246065, 0.1168440, 0.0093341, -0.0389239, -0.2061330, -0.1838580, -0.1319820, -0.2405010, -0.1042940, -0.0496872, -0.0359772, -0.1210220, -0.0432633, 0.0105878, 0.0031947, -0.0064133, 0.0000852, -0.0004026, 0.0027570, 0.0588290, 0.0577854, 0.0000611, 0.0042501, 0.0337514, 0.0509300, 0.0462826, 0.1874100, 0.2075390, 0.1886770, 0.2655690, 0.2836600, 0.1815290, 0.2774230, 0.3470130, 0.2295100, -0.0086284, -0.0343854, 0.1275740, -0.0184703, -0.1196700, -0.0783795, -0.0190984, -0.0231110, -0.0122729, -0.0002190, 0.0014564, 0.0123319, 0.0717766, 0.0498824, -0.0392578, 0.0646336, 0.0708016, 0.1242940, 0.1325020, 0.0952418, 0.1455050, 0.1837990, 0.1078990, 0.0647033, 0.1048940, 0.1906560, 0.1876920, 0.2272360, 0.1379690, 0.0224436, -0.0162374, -0.1109080, -0.0230116, -0.0497544, -0.0606983, -0.0421808, -0.0022498, 0.0078553, 0.0073276, 0.0165329, 0.0474915, 0.0317707, -0.0036868, 0.0801462, 0.1409230, 0.3652080, 0.1793010, 0.1953280, 0.1067680, 0.0703727, -0.0224816, 0.0655890, 0.0365078, 0.0810958, 0.0274406, 0.1614450, 0.0441120, -0.1207520, -0.2318110, -0.1026500, 0.0515063, -0.0565192, -0.1338180, -0.0171818, -0.0005859, 0.0002210, 0.0083365, 0.0250601, 0.0522558, 0.0558721, 0.0342042, 0.1734120, 0.2192110, 0.2208400, 0.0846437, 0.1847320, 0.1628720, 0.0845766, 0.0572732, 0.0647410, 0.0374460, -0.0209372, 0.0407971, 0.0270405, -0.0802797, -0.1992390, -0.1709310, 0.1198300, 0.1437410, 0.0530066, -0.0453798, 0.0089202, 0.0195264, 0.0003235, 0.0063255, 0.0494708, 0.0559311, 0.0601487, 0.1170900, 0.2816250, 0.2105820, 0.0617164, -0.0162010, -0.0583461, 0.1406190, -0.0853221, 0.1004750, 0.1655470, 0.2175800, 0.2430690, -0.0062536, -0.1310510, -0.1819730, -0.0773671, 0.1706260, 0.3834080, 0.2808920, 0.1082470, 0.0276547, 0.0165106, 0.0051871, 0.0001001, 0.0113054, 0.0521722, 0.0600286, 0.0955813, 0.0428011, 0.1750770, 0.1203880, -0.0273791, -0.2869500, -0.1908980, -0.0117633, 0.0324998, 0.1897120, 0.1472490, 0.1370260, 0.0141812, 0.0734346, -0.0736433, 0.0355485, 0.3541640, 0.4021380, 0.4475850, 0.3460980, 0.2049280, 0.0607888, 0.0061993, 0.0008461, 0.0000784, 0.0055488, 0.0380850, 0.0560647, 0.1232490, -0.0301336, 0.0672314, 0.0117135, 0.0723018, 0.0199622, -0.1757790, -0.0645007, 0.0024083, -0.1015310, -0.1104560, -0.0515437, -0.1141380, 0.0862934, 0.1419110, 0.3471340, 0.3487450, 0.2999920, 0.2094140, 0.2308610, 0.1389580, 0.0683341, 0.0111481, 0.0036438, -0.0003193, 0.0039562, 0.0199737, 0.0447394, 0.1145720, 0.0218243, 0.0835385, -0.0346196, -0.0273093, -0.0125641, 0.0128734, 0.0129509, -0.0162885, -0.1560920, -0.3044450, -0.3058510, -0.1930790, 0.1249530, 0.2016970, 0.2381790, 0.1109900, 0.1189310, 0.0623278, -0.0228496, 0.0912847, 0.0456483, 0.0163667, 0.0051617, -0.0001241, 0.0016793, 0.0096789, 0.0039019, -0.0112510, -0.0904399, 0.0224325, -0.0886878, -0.0422550, 0.0540540, 0.1286420, -0.0556608, -0.0812141, -0.2622820, -0.4763860, -0.2107510, -0.2660830, 0.0349016, 0.1798010, 0.1563030, 0.1273840, 0.0151030, -0.0036925, 0.0802053, 0.1138720, 0.0606363, 0.0365536, 0.0008863, 0.0000708, -0.0012949, -0.0009938, -0.0174046, -0.0597241, 0.0543808, -0.0114656, -0.0809012, -0.0082715, 0.1031220, 0.0785472, -0.0017103, -0.2155630, -0.3814980, -0.2380930, 0.1262970, -0.1151370, 0.1066000, 0.1648820, 0.0892374, 0.2146730, 0.0670690, -0.0182847, 0.1018040, 0.1677150, 0.0248071, -0.0144432, 0.0050445, -0.0004301, -0.0002788, 0.0020202, -0.0424232, 0.0303826, 0.0244070, -0.0663572, -0.0944141, -0.0403728, 0.0304406, 0.0623375, -0.0716437, -0.2366860, -0.2980430, -0.0997575, 0.1121160, 0.1135070, 0.1403320, -0.0567373, -0.0271228, 0.1729720, 0.0995163, 0.1276850, 0.0299577, 0.0056049, -0.0001197, 0.0369547, 0.0134178, -0.0003912, -0.0000772, -0.0149292, -0.0729081, -0.0034917, 0.0286434, -0.1064470, -0.2572520, -0.2610770, -0.1806220, 0.0101761, -0.0076644, -0.0252077, -0.1417430, -0.0854088, 0.2097420, 0.0369128, 0.0854974, -0.0510364, -0.0205938, 0.0785017, -0.0134510, 0.1234270, 0.0155143, 0.1262240, 0.0387630, 0.0226276, 0.0214155, 0.0015279, -0.0003939, -0.0124216, -0.1228910, -0.0703408, -0.0754620, -0.1877060, -0.1299800, -0.0780655, -0.2687960, -0.0359209, 0.0532133, -0.1190400, -0.2587950, -0.0361497, 0.0241305, 0.0491534, 0.0526000, 0.0391290, -0.0107989, -0.0796782, -0.0178352, 0.1837100, 0.0524152, 0.0984347, 0.0207318, 0.0128929, -0.0002765, 0.0005457, 0.0065908, -0.0016837, -0.1128220, -0.0926617, -0.1183710, -0.1528950, 0.0068570, 0.0248202, -0.1882250, -0.0251330, -0.0340450, 0.1865410, 0.0056857, -0.1202140, -0.1354850, -0.2854650, -0.0363547, -0.0112623, -0.0502954, -0.1214940, -0.0560952, 0.0906589, 0.0733091, 0.0483415, -0.0048428, 0.0019426, -0.0000236, 0.0004243, 0.0024054, -0.0013545, -0.0351762, -0.0114623, 0.1007640, -0.0312121, -0.0095435, 0.0446173, -0.0765171, 0.1268670, 0.0797868, 0.0946452, -0.0160807, -0.3777880, -0.2859430, -0.4205570, -0.1223010, -0.1728740, -0.1818050, -0.2701230, -0.1654750, -0.0862873, 0.0069694, 0.0503253, 0.0228896, -0.0014401, -0.0004589, 0.0004142, -0.0001201, -0.0011416, -0.0138846, -0.0292315, 0.0739137, 0.1113330, 0.0874092, -0.0354654, 0.0916059, 0.0895856, 0.0273332, -0.0190265, -0.1475760, -0.2479600, -0.1975590, -0.1791380, -0.1902140, -0.2808420, -0.3680120, -0.3929150, -0.3221580, -0.1549850, -0.0161029, 0.0130820, 0.0219464, 0.0066419, 0.0001936, 0.0001025, 0.0005475, 0.0001436, -0.0016768, -0.0345074, 0.0119919, 0.1408940, 0.2433880, 0.2388350, 0.2417580, 0.1743600, 0.1020770, 0.2319950, 0.0921819, 0.1097410, 0.0258835, -0.0159508, -0.1287320, -0.1909580, -0.3212640, -0.3086500, -0.3630990, -0.0972400, -0.0084517, 0.0138458, 0.0150751, -0.0027303, -0.0007781, 0.0001860, 0.0001544, -0.0049112, -0.0185725, -0.0350778, 0.0336044, 0.1281410, 0.1860960, 0.1190200, 0.1364310, 0.1956600, 0.2391850, 0.1679400, 0.0804001, 0.1287630, 0.0325416, 0.0647793, 0.0631731, -0.1467930, -0.1805270, -0.1991680, -0.2190090, -0.0126346, 0.0300317, 0.0386626, 0.0019993, -0.0061113, -0.0000745, -0.0003263, 0.0000608, -0.0071267, -0.0115197, 0.0130743, 0.0673045, 0.0407013, 0.0506237, -0.0226858, -0.0747774, 0.0479541, -0.0653593, -0.0056590, 0.0144174, 0.0251179, -0.0173554, -0.0663694, -0.0631530, -0.0609504, 0.0375210, -0.0030105, -0.0524250, 0.0096328, 0.0440261, 0.0315350, 0.0014453, 0.0002764, -0.0004848, -0.0001824, 0.0001913, -0.0013286, 0.0049051, 0.0330260, 0.0457145, 0.0401912, 0.0426146, 0.0238416, -0.0299734, 0.0457065, 0.0418463, -0.0027081, -0.0705766, 0.0710109, 0.0633827, 0.0855331, 0.0311950, 0.0509364, 0.1689150, 0.0595197, 0.0253431, 0.0047361, 0.0103339, 0.0125116, -0.0001260, 0.0001733, -0.0000349, 0.0000924, -0.0002105, 0.0000471, 0.0004571, 0.0029913, 0.0131422, 0.0386191, 0.0508536, 0.0663286, 0.0693930, 0.0705977, 0.0648419, 0.0811195, 0.0832746, 0.0417295, -0.0120912, 0.0224942, 0.0265395, 0.0730286, 0.0867668, 0.0637085, 0.0503946, 0.0251976, 0.0039704, 0.0027983, 0.0000235, 0.0006154, 0.0000136, -0.0009333, -0.0000024, 0.0005299, -0.0002071, -0.0004865, -0.0004240, 0.0026066, 0.0152458, 0.0143674, 0.0031163, 0.0099673, 0.0034176, 0.0006210, 0.0039422, 0.0052551, -0.0022315, 0.0157155, 0.0219344, 0.0482149, 0.0193742, 0.0087337, 0.0189513, 0.0127178, 0.0001830, 0.0004771, 0.0001603, -0.0000100, -0.0003725, -0.0002368, -0.0000268, -0.0001871, -0.0001666, 0.0002458, -0.0000814, 0.0002621, 0.0004575, -0.0000095, 0.0000202, 0.0000876, -0.0004195, 0.0000809, 0.0001201, 0.0005263, 0.0003775, -0.0002802, -0.0002610, -0.0001168, -0.0003387, -0.0005674, -0.0000488, -0.0001144, 0.0007747, -0.0003114, 0.0003384, 0.0002984, 0.0002532, 0.0002414, -0.0005892, 0.0004316, -0.0003824, -0.0000190, 0.0002561, 0.0000299, -0.0005125, -0.0011947, -0.0023275, -0.0027501, -0.0029977, -0.0043754, 0.0009133, 0.0104609, 0.0078092, 0.0170517, 0.0049212, -0.0028332, -0.0040220, -0.0047818, -0.0033315, -0.0002217, -0.0005190, 0.0003664, -0.0006256, 0.0001881, 0.0000323, 0.0001911, 0.0006740, 0.0003702, 0.0003505, 0.0002494, -0.0001446, -0.0002275, -0.0015921, 0.0032829, 0.0323504, 0.0221693, -0.0247964, -0.0216425, 0.0337825, 0.0147958, 0.0499308, 0.0626104, -0.0011520, -0.0032037, -0.0407575, -0.0319758, -0.0437754, -0.0312967, -0.0132194, 0.0016077, 0.0052659, -0.0000279, -0.0004592, -0.0004005, -0.0007289, 0.0061161, 0.0024304, 0.0055008, -0.0037476, -0.0019920, -0.0109104, 0.0289988, 0.1034190, 0.1277140, 0.0186501, 0.0899616, 0.1292030, -0.0375817, 0.0383209, 0.1685770, 0.1573170, 0.0784664, -0.0181162, 0.0219946, -0.0499537, -0.1022780, -0.0461450, -0.0307242, -0.0049039, -0.0128880, 0.0003331, -0.0003970, -0.0004055, 0.0206299, 0.0043575, -0.0064982, -0.0044757, 0.0306958, 0.1068010, 0.1457290, 0.2339010, 0.2278320, 0.2600520, 0.2102790, 0.0212980, 0.1226490, 0.0607917, -0.0296742, 0.0081823, 0.0551192, -0.0116221, 0.0423208, 0.0396724, -0.0801657, -0.0032090, 0.0853747, 0.0050815, -0.0038994, -0.0091146, 0.0001224, 0.0000155, 0.0025976, 0.0053022, -0.0223029, 0.0015975, 0.0511937, 0.0801602, 0.0675149, 0.1609380, 0.2217710, 0.4483960, 0.3919510, 0.2431990, 0.1843490, 0.1225040, 0.3266220, 0.2867360, 0.1339520, 0.1373940, 0.3303710, 0.1622220, 0.1178750, 0.0135455, -0.0035542, 0.0003025, -0.0104720, -0.0137960, 0.0003702, -0.0003749, -0.0023461, -0.0053537, -0.0853768, -0.0654532, -0.0031804, 0.0419392, 0.0947477, 0.3021590, 0.4088180, 0.3465900, 0.4369600, 0.4150880, 0.5550050, 0.4620120, 0.4168610, 0.4536490, 0.3290770, 0.1721670, 0.2961630, 0.0330968, 0.0012038, 0.1117530, 0.0479821, -0.0207316, 0.0138762, -0.0110476, 0.0003965, -0.0032491, -0.0087597, -0.0374328, -0.1143040, -0.0604369, -0.0385348, 0.0184039, 0.2295000, 0.1736350, 0.1799350, 0.1781520, 0.2140810, 0.0519382, 0.1476340, 0.0351968, 0.2117200, 0.0744233, 0.0302126, -0.1341670, -0.0538823, -0.0964025, -0.0385880, -0.0014389, -0.0038130, 0.0636043, 0.0100676, -0.0058094, -0.0013345, -0.0049441, -0.0184336, -0.0435393, -0.1019570, -0.0883306, 0.0266007, 0.0575124, 0.2814330, 0.0166262, -0.0833432, -0.0563177, -0.2000380, -0.2412000, -0.2720430, -0.2670480, -0.3008520, -0.2687920, -0.1089500, -0.0452289, -0.3499380, -0.1118650, 0.0023232, 0.1571900, 0.2135130, 0.1477310, 0.0297937, 0.0031509, 0.0000173, -0.0080496, -0.0169391, -0.0256915, -0.0877049, -0.0726682, 0.0655247, 0.0312873, 0.1450320, -0.0454955, -0.2398300, -0.1221000, -0.2602520, -0.3897960, -0.2755860, -0.0779834, -0.1066680, -0.1215770, 0.1133380, 0.1544260, -0.1471430, 0.0176329, 0.1468460, 0.0920115, 0.1060910, 0.1288730, 0.0689418, -0.0008259, -0.0000343, -0.0055015, -0.0209115, -0.0320415, 0.0508442, 0.0659482, 0.0978591, 0.0232958, 0.0068750, -0.2292040, -0.2747170, -0.0983099, 0.0565726, -0.1881760, -0.0749101, 0.0060442, 0.1802770, 0.0740050, 0.2137390, 0.2251900, -0.0418613, 0.0787741, 0.1131210, 0.0896883, 0.0360256, 0.1171530, 0.0456821, -0.0016933, -0.0006234, -0.0063507, -0.0416057, -0.0645077, 0.1091220, 0.0588521, 0.0676951, -0.0887543, -0.4106150, -0.4825370, -0.3727630, -0.2000150, 0.1242030, -0.2257540, 0.0420606, 0.2809360, 0.3073570, 0.2134850, 0.1393750, 0.1513670, -0.0728623, -0.0910447, -0.0849949, -0.0002579, 0.0421620, 0.0863060, 0.0302740, -0.0003556, -0.0002308, -0.0041861, -0.0389873, -0.0180265, 0.1378630, -0.0136882, -0.0704717, -0.2319850, -0.5443710, -0.3533970, -0.0680068, -0.0072117, -0.0674104, -0.0269618, 0.2781660, 0.2904260, 0.0562441, 0.0253207, -0.0817665, 0.0968470, -0.0028570, -0.0629902, -0.2331690, -0.2880220, -0.2361360, -0.0504725, 0.0050701, -0.0007874, -0.0002653, -0.0017450, -0.0272432, 0.0061106, 0.0372927, 0.0354653, -0.1478500, 0.1108090, -0.1796710, -0.2771110, -0.3962610, -0.0472367, 0.0139057, 0.1161850, 0.1707660, 0.0531134, 0.1217930, 0.1582600, -0.0110370, -0.0315697, 0.0888370, -0.0123343, -0.1419720, -0.3576630, -0.2550830, -0.0581130, 0.0040371, 0.0006197, -0.0004888, -0.0015874, -0.0134264, 0.0137901, 0.0431566, -0.1446040, 0.0444710, -0.0427461, -0.1845580, -0.3337390, -0.3085010, -0.1956670, -0.2048090, 0.1023860, 0.2391470, 0.0485673, 0.1124830, -0.0498527, 0.0816222, -0.2584830, -0.2106500, -0.2156500, -0.2007980, -0.2936940, -0.2190350, -0.0506291, 0.0109970, 0.0002780, -0.0003487, 0.0000031, 0.0020602, 0.0134078, 0.0572979, -0.1381490, -0.0703592, -0.2565600, -0.2468400, -0.2034680, -0.2892650, -0.1996450, -0.2212200, 0.1331730, 0.0661087, 0.0437284, 0.0262721, -0.2309910, -0.1321930, -0.2274950, -0.3508670, -0.2646190, -0.2820680, -0.2096480, -0.1859800, -0.0260637, 0.0163687, 0.0053795, 0.0004865, -0.0000900, 0.0059792, 0.0133135, 0.0258477, -0.0015508, 0.0839337, -0.2182590, -0.2422670, -0.0900715, -0.2436640, -0.5085900, -0.0750324, 0.1035030, 0.1286370, 0.0560560, -0.0933105, -0.0625352, -0.1129230, -0.1770880, -0.1668000, -0.0612826, -0.0463799, -0.0606751, -0.0856295, 0.0326092, 0.0425383, 0.0154349, -0.0002422, 0.0002196, 0.0040015, 0.0948192, 0.1807500, 0.1639370, 0.2369020, -0.2194950, -0.0232848, -0.0413732, -0.2804450, -0.4960130, -0.2859180, -0.1625440, 0.0864556, 0.1955580, -0.1589110, 0.0821932, 0.0553405, -0.0455133, -0.0321313, -0.0241501, -0.1476980, -0.0551458, -0.0489397, 0.0337554, 0.0174285, 0.0069281, -0.0007763, 0.0001717, 0.0002793, 0.1076510, 0.2247950, 0.3169870, 0.3763640, -0.0787482, -0.2301400, -0.1851570, -0.0508929, 0.0407247, -0.3112020, -0.2293410, 0.1106660, -0.0877309, -0.0229147, 0.0906486, -0.0939281, 0.1101100, 0.1414930, 0.0294632, -0.0003463, 0.1236630, 0.1708360, 0.0504181, -0.0039024, 0.0036202, -0.0003313, -0.0005719, 0.0061314, 0.0299120, 0.1307320, 0.2322550, 0.3358350, 0.2346460, 0.1501340, 0.1572430, 0.1220550, 0.0819031, 0.0012432, 0.0623775, -0.0557652, 0.1309020, 0.2304140, 0.0519724, -0.0511990, 0.1399770, 0.0287166, -0.0392834, 0.0291772, 0.2432650, 0.2285820, 0.0564011, 0.0108903, -0.0000066, 0.0006325, -0.0012761, 0.0083655, 0.0235461, 0.0954110, 0.2214190, 0.3626470, 0.1949210, 0.4091540, 0.1153090, 0.1289110, 0.1480470, 0.0317087, 0.0558188, -0.2921430, -0.0757726, 0.2703520, 0.0548119, 0.0951519, 0.1181350, -0.0437129, -0.0347931, 0.1913870, 0.2053380, 0.1276590, 0.0296915, 0.0022392, -0.0002050, 0.0004547, -0.0005893, 0.0096239, 0.0136306, 0.0715526, 0.1510670, 0.1431640, 0.1814400, 0.1137380, 0.1570050, 0.1035150, -0.0611422, -0.1957050, -0.1145900, -0.2781510, -0.1443420, 0.0791093, 0.0444810, 0.1687980, 0.2607710, 0.2119170, 0.2837760, 0.1881560, 0.1875110, 0.1193660, 0.0661144, 0.0049494, 0.0004259, 0.0000622, -0.0006186, -0.0005458, 0.0162972, 0.0418979, -0.0027875, 0.0242466, 0.0716220, 0.0519273, 0.0505981, -0.0177769, -0.0254807, -0.0592091, -0.1897630, 0.0448484, -0.0007038, -0.1014330, 0.1687930, 0.2134740, 0.0803993, 0.2373780, 0.1146610, 0.0885422, 0.1919940, 0.1336660, 0.0733908, 0.0202653, -0.0003581, 0.0001911, 0.0003204, 0.0034067, 0.0147653, -0.0146542, -0.0727337, -0.1540580, -0.1089620, 0.1452080, 0.0576679, -0.0524233, -0.0599376, 0.0237922, 0.0345968, -0.0563322, 0.1616870, 0.2066830, 0.1239570, -0.0072144, 0.0802450, 0.1593280, 0.0531174, 0.1104410, 0.1500840, 0.0935407, 0.0633599, 0.0122814, -0.0002849, 0.0000731, 0.0000476, 0.0078421, 0.0047007, -0.0573866, -0.1223820, -0.1243870, -0.0189380, 0.0428779, -0.0728400, -0.0421453, -0.0986234, -0.0987039, -0.1050860, -0.2293610, -0.0123595, 0.1215070, -0.0289407, 0.0761808, 0.0535859, 0.0036543, -0.0172944, 0.0320113, 0.0408416, 0.0127314, 0.0003371, -0.0000795, 0.0001664, 0.0001032, -0.0000276, 0.0021358, -0.0071604, -0.0428288, -0.0896620, -0.1106830, -0.1255160, -0.0668073, -0.1188830, -0.1041020, -0.1058730, -0.0202405, -0.0103759, 0.0246444, -0.0364910, -0.0055217, -0.0166517, 0.0036711, 0.0489803, 0.0554174, 0.0413607, -0.0020004, -0.0077215, 0.0031691, 0.0002209, 0.0000022, 0.0001884, -0.0003208, 0.0001249, 0.0001900, -0.0001596, 0.0010420, -0.0093013, -0.0112987, -0.0028485, 0.0087918, 0.0196948, 0.0311093, 0.0166333, -0.0012251, -0.0435316, -0.0647699, -0.0714657, -0.0564540, -0.0526647, -0.0584032, -0.0316352, 0.0011541, 0.0451345, 0.0054522, 0.0008680, 0.0000588, -0.0005271, 0.0002625, 0.0003000, 0.0001949, 0.0001891, -0.0004121, 0.0003633, -0.0000983, -0.0006196, 0.0000098, -0.0008689, -0.0007787, -0.0008620, -0.0123458, -0.0034608, -0.0021397, -0.0036882, -0.0050453, -0.0079586, -0.0151993, -0.0119135, -0.0043280, -0.0081729, -0.0050487, 0.0009412, 0.0046518, 0.0003638, 0.0002978, -0.0002655, 0.0003413, 0.0000746, 0.0000864, 0.0001895, 0.0000064, 0.0003255, 0.0005839, -0.0004540, -0.0004084, -0.0003365, -0.0007639, -0.0002985, -0.0002833, 0.0004910, 0.0000910, 0.0001318, -0.0005568, -0.0004193, -0.0000952, -0.0002073, 0.0001291, -0.0001529, -0.0007060, -0.0000889, 0.0001398, -0.0000465, 0.0001813, 0.0001148, 0.0001515, 0.0001420, 0.0001335, -0.0004401, -0.0001578, -0.0005425, -0.0002734, 0.0000299, 0.0002236, 0.0000282, 0.0011393, 0.0007217, 0.0007536, -0.0007566, -0.0016496, 0.0057886, -0.0055298, -0.0131722, 0.0255715, 0.0046022, -0.0029477, -0.0081094, -0.0159156, -0.0144743, -0.0019589, 0.0000389, 0.0001627, -0.0000273, -0.0000015, 0.0002848, 0.0006979, 0.0001260, 0.0000801, 0.0007130, 0.0002159, 0.0006520, -0.0005000, -0.0004516, 0.0096416, 0.0259100, 0.0292354, 0.0167459, 0.0191575, -0.0002480, -0.0075820, -0.0764627, -0.0814070, -0.0542916, -0.0459762, -0.0664055, -0.0661090, -0.0664289, -0.0356058, -0.0099550, 0.0029305, 0.0047179, 0.0005221, 0.0010545, 0.0001352, -0.0002469, 0.0004514, 0.0019047, 0.0005313, 0.0053042, 0.0045845, 0.0105832, 0.0594537, 0.0898694, 0.1553240, 0.1891700, 0.2075180, 0.1195200, -0.0130930, 0.0219866, 0.1873870, 0.0947894, -0.0421966, -0.0881001, -0.0443558, -0.1425670, -0.1547100, -0.0890259, -0.0332645, 0.0071205, 0.0013406, -0.0002450, 0.0002788, 0.0001512, 0.0028504, 0.0022961, 0.0029862, 0.0206404, 0.0504172, 0.1305070, 0.2623470, 0.2735360, 0.3305550, 0.3262660, 0.3258440, 0.2119000, 0.1902780, 0.3429970, 0.2028740, 0.0024201, -0.0246008, -0.0717773, -0.1067000, -0.2026080, -0.2138720, -0.1875410, -0.0185569, 0.0186857, 0.0098377, -0.0049113, 0.0005800, -0.0004975, 0.0009330, 0.0057270, 0.0147883, 0.0251326, 0.1004120, 0.2046650, 0.3063300, 0.4345570, 0.5402310, 0.2820860, -0.0254491, -0.0386550, -0.0451402, 0.0510810, 0.1417470, -0.0045343, 0.1195060, 0.0907017, -0.0010022, -0.1369570, -0.1253920, -0.2025990, -0.0822652, -0.0149110, -0.0051016, -0.0090146, -0.0000576, -0.0001714, 0.0070684, 0.0168565, 0.0017087, -0.0209372, 0.1627990, 0.3531700, 0.4446090, 0.5161710, 0.3318970, 0.0074062, -0.1948840, -0.1786990, -0.2375030, -0.0436005, 0.1277240, 0.0989963, 0.0957509, 0.0865756, -0.0114744, -0.0465543, -0.0926173, -0.1511130, -0.0485603, 0.0155641, 0.0214930, -0.0010992, -0.0004343, 0.0053286, 0.0207920, 0.0265181, 0.0285837, 0.0147467, 0.1896670, 0.3671870, 0.6270140, 0.3670180, 0.0670450, -0.1429400, -0.2306720, -0.2691110, -0.1394120, 0.2067540, 0.3496140, 0.0373329, 0.0730132, 0.0542569, 0.0906207, 0.1690320, -0.1106380, -0.1915520, -0.0589146, 0.0173640, -0.0231472, 0.0002058, -0.0006073, -0.0010502, 0.0168230, 0.0244276, 0.0492150, 0.0221763, 0.0091943, 0.0799766, 0.3793970, 0.5102960, 0.3568800, -0.1708870, -0.4708310, -0.2806290, -0.1482670, 0.2094040, 0.4150900, 0.1920400, 0.2227480, 0.1352010, 0.2148810, 0.1002780, -0.0163107, -0.0367287, -0.1429210, -0.0853967, -0.0157522, 0.0028498, 0.0002326, -0.0000322, 0.0081943, 0.0392441, 0.0765586, 0.0385971, 0.0277933, 0.0908360, 0.3668150, 0.4860970, 0.2895360, -0.0953143, -0.2630180, -0.1584460, -0.2038800, -0.0656038, 0.1372960, 0.2892490, 0.1878210, 0.2942670, 0.3232030, -0.0086712, 0.0818008, 0.0116619, -0.1088070, -0.0134743, 0.0252304, -0.0011541, -0.0001552, 0.0003374, 0.0052231, 0.0423827, 0.0866103, 0.1387100, 0.0486670, 0.1813740, 0.2351110, 0.1909310, 0.1718130, 0.0751268, -0.0901276, -0.1382920, -0.2703880, -0.2794500, 0.2301650, 0.1447410, 0.0959703, 0.0947924, 0.1368480, 0.0519871, 0.0889593, 0.1264750, 0.0266377, 0.0216458, 0.0493657, -0.0008108, 0.0003044, 0.0009721, -0.0016829, 0.0294843, 0.0670560, 0.1076670, 0.0879723, 0.1581720, 0.1368290, -0.0588836, -0.2675850, -0.0803559, -0.2398000, -0.0227408, -0.1067100, -0.2107790, -0.0132157, 0.2781320, 0.0898801, 0.0174871, 0.0478409, 0.0093713, 0.0999165, 0.0696441, 0.0859789, 0.0928453, 0.0301552, 0.0004336, -0.0002326, 0.0004170, -0.0039724, 0.0100460, 0.0662090, 0.1126420, 0.1839490, 0.1491130, 0.0352303, 0.0828101, 0.0492848, -0.4355580, -0.4887460, -0.3014960, -0.0412738, -0.2110460, 0.0753670, 0.1716380, 0.1892980, 0.1436980, -0.2019250, -0.2024330, -0.0010697, 0.0151519, 0.0383865, 0.1012770, 0.0489281, 0.0019884, -0.0001373, 0.0005561, -0.0036122, 0.0192208, 0.0879419, 0.1408670, 0.2101700, 0.0194897, 0.0110410, -0.0146363, 0.1231670, -0.2313030, -0.4561630, -0.0856781, -0.1072310, -0.3545910, -0.0321666, 0.1155730, 0.1049310, 0.0674947, -0.2124240, -0.0738732, 0.0626245, 0.0936675, 0.1393740, 0.0980459, 0.0789839, 0.0125775, -0.0006840, 0.0021072, 0.0003352, 0.0188175, 0.0529775, 0.1159440, 0.2434370, 0.0719218, -0.0194171, 0.1160280, 0.0039149, -0.0986768, -0.1506320, 0.0107864, -0.1814350, -0.1859700, 0.0450670, 0.2272260, 0.1404320, 0.0278656, -0.0414326, -0.0662630, 0.1004860, 0.2454240, 0.2303780, 0.0929828, 0.0834718, 0.0004483, -0.0003311, 0.0036332, 0.0038037, 0.0003753, 0.0019806, 0.1077910, 0.0677147, 0.0416102, 0.0310135, 0.2247670, 0.0997716, -0.0231950, 0.0429480, -0.0807187, -0.5243210, -0.2547050, 0.1303020, 0.1657510, 0.0377716, 0.0791255, 0.1240600, -0.0842459, 0.0840415, 0.1952420, 0.2460220, 0.1421560, 0.0636908, 0.0102322, -0.0005527, 0.0013390, 0.0095191, 0.0017924, -0.0097375, 0.0004542, 0.0748537, 0.0838463, -0.0461558, 0.1017720, -0.0144261, -0.1413400, 0.0206794, -0.1569580, -0.2533150, -0.1003460, 0.0498942, 0.1556320, 0.0834946, 0.0360963, 0.2345090, 0.1823360, 0.2424640, 0.2493200, 0.1797660, 0.1715270, 0.1169760, 0.0249831, 0.0003838, 0.0004924, 0.0105931, 0.0112197, -0.0175432, 0.0080538, 0.0074781, -0.0041847, -0.0964931, -0.0714777, -0.2235260, -0.0441811, 0.0063638, -0.1194550, -0.0719264, 0.0107860, 0.2656280, 0.1629160, 0.0489492, 0.0826975, 0.1144500, 0.0572567, 0.1584960, 0.1317480, 0.1064400, 0.1127250, 0.0565640, 0.0207063, 0.0011165, 0.0001134, 0.0099312, 0.0463332, -0.0173212, 0.0312558, 0.0615871, -0.1315990, 0.0167683, -0.1741840, 0.0109862, 0.0445151, -0.1582250, -0.1559240, -0.0040884, 0.0458309, 0.0311767, 0.0927545, 0.0665527, -0.0456246, 0.0000989, 0.1046740, 0.2600150, 0.1626480, 0.1059580, 0.0176319, -0.0063362, 0.0031075, -0.0000996, 0.0016662, 0.0023365, 0.0745356, 0.1111870, 0.0502121, 0.0058915, -0.0005645, 0.0265040, -0.0757467, -0.0741853, -0.2122640, -0.1438830, 0.0917821, 0.0727391, 0.0278086, 0.0297945, 0.2228280, 0.2250010, 0.0535830, -0.0070538, 0.1024500, 0.2475930, 0.1636430, 0.0333515, -0.0064058, 0.0156283, -0.0003553, -0.0001034, -0.0010220, 0.0015962, 0.1029680, 0.2497060, 0.0675678, -0.0778407, 0.0722696, 0.0856396, 0.0615324, -0.0677994, -0.1938940, -0.1466340, 0.1700680, 0.0401303, -0.0242606, 0.1146920, 0.0536400, 0.0357649, -0.0362910, 0.0900554, 0.2043520, 0.2106120, 0.0891072, -0.0001048, -0.0141419, 0.0047879, 0.0003752, 0.0002821, 0.0008058, 0.0071837, 0.0703916, 0.1822640, 0.0341516, -0.0785693, 0.1192460, -0.1210170, -0.2287960, -0.0138689, -0.1163410, -0.1237860, -0.0489935, 0.1086430, 0.2554980, 0.2469630, 0.0470563, 0.0466135, 0.1103110, 0.1467040, 0.1906190, 0.1756670, 0.0628075, -0.0169003, 0.0088479, 0.0002749, -0.0001450, 0.0000605, 0.0007169, 0.0053101, -0.0111228, 0.0337336, 0.0017768, 0.1017250, 0.0606406, -0.0671847, -0.0075864, -0.0091836, -0.0783661, -0.1600230, -0.1410890, 0.0198526, 0.1639510, 0.0160107, -0.0474193, 0.0698349, 0.0078269, 0.0427801, 0.0722107, 0.1107430, 0.0354609, 0.0048889, 0.0006252, -0.0000981, 0.0003479, -0.0001847, -0.0002822, 0.0066164, 0.0571468, 0.0310728, -0.0380460, -0.0722513, -0.0387837, -0.0853204, 0.0030765, 0.0689764, -0.1360240, -0.2998130, -0.1689900, -0.1804280, 0.0554365, 0.0959339, 0.1753320, 0.0443426, -0.0871907, -0.0521362, 0.0289227, 0.0728111, 0.0300197, 0.0109532, -0.0023057, -0.0005915, 0.0001555, -0.0004936, -0.0000915, 0.0020210, 0.0402851, 0.0521701, -0.0147755, 0.0483337, -0.0050426, 0.0506216, -0.0094711, 0.0728871, 0.0052952, 0.0123952, -0.0662422, 0.0050843, 0.0075042, 0.1038340, 0.2055070, 0.0128746, -0.0554760, -0.0807426, 0.0181035, -0.0090352, -0.0146304, -0.0014102, -0.0033441, -0.0001882, -0.0000501, -0.0000466, -0.0001163, -0.0002463, -0.0123736, -0.0264065, 0.0106535, 0.0671485, 0.0855810, 0.1766220, 0.0936772, 0.0009711, -0.0147695, 0.1796610, 0.0558376, 0.0861827, 0.1598210, 0.2701090, 0.2538550, 0.1440790, 0.0925673, -0.0376109, -0.0387361, -0.0543071, -0.0431727, -0.0025954, -0.0007187, -0.0005759, -0.0004017, 0.0001957, 0.0002678, -0.0000071, -0.0001114, 0.0043203, 0.0023875, 0.0126461, 0.0465237, 0.0524030, 0.0412746, 0.0805856, 0.0923002, 0.0820507, 0.1080510, 0.1108740, 0.0916156, 0.0883391, 0.1084730, 0.0963230, 0.0386798, 0.0392952, 0.0132551, 0.0015668, -0.0001720, -0.0001799, 0.0001534, 0.0004979, -0.0000367, 0.0001006, 0.0001614, 0.0001469, 0.0000974, -0.0002383, -0.0005629, 0.0012146, 0.0090396, 0.0082715, 0.0026168, 0.0017735, 0.0042591, 0.0080241, 0.0046107, 0.0225867, 0.0028926, 0.0011562, 0.0058359, 0.0191032, -0.0015568, -0.0007952, 0.0002593, -0.0000540, -0.0001085, 0.0001016, 0.0000627, 0.0001517, -0.0000676, 0.0002461, 0.0002595, 0.0003255, 0.0001302, -0.0005557, -0.0000233, -0.0002114, 0.0005813, -0.0002499, -0.0000478, -0.0003094, -0.0001018, -0.0001471, -0.0007896, 0.0004140, -0.0000253, 0.0003373, -0.0003624, 0.0004645, -0.0000514, 0.0001573, 0.0003370, 0.0001580, -0.0000472, -0.0002135, 0.0000630, -0.0000611, -0.0000895, 0.0005140, -0.0001147, 0.0007375, -0.0007178, -0.0000588, -0.0004006, -0.0006755, -0.0008964, -0.0015764, -0.0008629, -0.0029149, 0.0005479, -0.0047354, -0.0045236, -0.0003162, -0.0131893, -0.0119075, -0.0109424, -0.0124839, -0.0099722, -0.0093251, -0.0075797, -0.0007286, 0.0002170, 0.0001391, -0.0001122, -0.0000359, -0.0006677, 0.0000763, -0.0006358, 0.0006154, -0.0017212, -0.0007278, -0.0000198, 0.0010649, 0.0028999, 0.0130944, 0.0427688, 0.0513848, 0.0460732, 0.0702480, 0.0795927, 0.0503969, -0.0238516, -0.0333265, -0.0038833, -0.0030261, -0.0301592, 0.0071490, 0.0074347, 0.0019287, -0.0003686, 0.0043653, 0.0027359, 0.0000750, -0.0001883, 0.0003441, -0.0003187, -0.0004104, -0.0053553, -0.0082629, -0.0193489, -0.0124810, -0.0106129, -0.0071705, 0.0594786, 0.0013401, -0.0283069, -0.0549395, 0.0557569, 0.0389907, -0.0119195, 0.0142276, -0.0738573, -0.0800511, -0.0064154, -0.1209770, 0.0183062, 0.0586640, 0.0481153, 0.0118709, -0.0064354, -0.0041681, 0.0002679, -0.0006009, 0.0004989, 0.0000705, -0.0007380, 0.0003830, -0.0210332, 0.0255031, 0.0325024, 0.0071514, 0.0023600, -0.0430952, -0.1403360, -0.0623823, -0.0468931, 0.2171800, 0.1993000, 0.1579130, 0.0590224, -0.0798346, -0.0114626, -0.0406738, 0.1083400, 0.1069350, 0.0368646, 0.0013783, 0.0039726, 0.0074107, 0.0014638, -0.0000462, -0.0004191, 0.0002568, -0.0080100, 0.0036041, 0.0151525, 0.0396162, 0.0406373, 0.0811975, 0.0081971, -0.0210573, 0.0083984, 0.2723260, 0.1361870, 0.0526932, -0.1648010, -0.0211661, 0.0134994, -0.0949157, -0.0332419, 0.0660601, 0.0960338, 0.0350293, -0.0255850, -0.0206504, 0.0237744, 0.0029218, 0.0012215, -0.0001973, -0.0000605, 0.0007334, 0.0146633, 0.0030374, 0.0376056, 0.0885826, 0.1404220, 0.0886578, 0.0880476, 0.1459840, 0.1785790, 0.1700540, 0.0512483, 0.0257938, 0.2044890, 0.0895055, -0.0152975, -0.0876624, 0.0146996, 0.0678085, 0.1309810, -0.0316776, -0.0303437, -0.1497810, -0.0268268, -0.0400982, -0.0005473, 0.0000595, -0.0022045, 0.0033746, -0.0062656, 0.0159566, 0.0631534, 0.1559100, 0.1689280, 0.1354310, 0.1757840, 0.1390720, 0.0653197, 0.1476570, 0.2864210, 0.0337257, -0.0457890, -0.0042363, 0.0026711, -0.0447522, -0.0014805, 0.0770582, 0.2268370, 0.0455221, -0.0799497, -0.0559885, -0.0001786, -0.0570708, -0.0035176, -0.0092683, 0.0031295, 0.0179108, 0.0019430, 0.0482517, 0.0818488, 0.1721570, 0.1992410, 0.1657230, 0.2178420, 0.0895038, 0.1248240, 0.1303790, 0.1446570, -0.1215240, -0.1150380, 0.0088205, 0.0416685, 0.0250449, 0.1647570, -0.0404321, -0.1457560, -0.0378441, 0.0608701, -0.1110220, -0.0753535, -0.0292288, -0.0043193, 0.0004038, 0.0018637, 0.0069170, 0.0053388, -0.0025587, 0.0737597, 0.1159720, 0.0553260, 0.0279247, 0.2239150, 0.1024420, 0.1401480, 0.1891520, 0.0536775, 0.0162752, -0.0293385, -0.0781360, 0.0246275, 0.0408444, -0.0380838, -0.0679193, -0.1234340, -0.0446407, -0.0327333, -0.0869480, -0.0843246, -0.0150848, -0.0020086, -0.0003906, 0.0009222, -0.0068548, -0.0538790, -0.0907946, 0.0308169, 0.0650820, -0.0964516, 0.0642994, 0.0431541, -0.0549220, -0.0392327, -0.0835853, -0.1702320, -0.1673280, -0.3400270, -0.3180470, -0.2379590, 0.1406600, 0.1059470, 0.0050393, -0.0761338, 0.0051828, 0.0293317, 0.0211558, -0.0967086, -0.0153689, 0.0018276, 0.0002037, 0.0013722, 0.0120862, -0.0553796, -0.0529982, 0.0056641, -0.0224178, -0.0751355, -0.0104272, 0.2274090, 0.1149800, -0.0880404, -0.0317676, -0.2154780, -0.1248930, -0.1449730, -0.0311079, -0.1936110, 0.1268240, 0.0323156, 0.2107380, 0.0207092, 0.1002290, 0.2155180, 0.1722630, 0.0405317, 0.0239158, -0.0008847, -0.0002436, 0.0002770, 0.0114836, 0.0065130, -0.0008943, 0.0070146, 0.0399820, -0.0053298, -0.0260516, 0.1464900, -0.0252236, -0.1950940, -0.3845500, -0.3016680, -0.3036750, -0.0964694, -0.0873010, 0.0917657, 0.0235139, 0.0362569, 0.2428380, 0.2106820, 0.0101325, 0.1814880, 0.1367980, 0.0555527, -0.0061269, 0.0004363, 0.0005075, 0.0006979, 0.0101625, -0.0277479, -0.0057836, -0.0458761, -0.0665748, -0.0894714, -0.0156716, 0.0887150, -0.0809464, -0.1787310, -0.3142950, -0.1133850, 0.0190707, 0.1006910, -0.0797212, 0.0435845, -0.0986053, -0.0419023, 0.1463960, 0.1273040, 0.0743309, 0.0949746, 0.0829079, 0.0543356, 0.0198593, 0.0084041, 0.0000997, 0.0003832, 0.0030415, -0.0218224, 0.0032493, -0.1162920, -0.0538414, 0.0929440, 0.0663455, -0.1577060, -0.0538290, -0.1056140, -0.2689340, -0.0288227, 0.2580960, 0.0650110, 0.1057600, 0.0674385, 0.1077830, -0.0628228, -0.1192940, 0.0133063, -0.0666261, 0.0550711, 0.0272298, 0.0904327, 0.0236723, 0.0000980, 0.0000873, -0.0001418, 0.0079899, 0.0118959, -0.0943293, -0.2073670, -0.0258158, 0.0506732, 0.0586665, -0.1226910, 0.0666647, 0.1273580, -0.2487670, 0.1798190, 0.3488410, 0.2146030, 0.1238200, -0.0678540, -0.1615700, -0.1903780, -0.2750900, -0.0454164, -0.1343130, -0.0518947, 0.0638107, 0.1109730, 0.0438236, 0.0048788, 0.0003832, -0.0002567, 0.0150870, -0.0267131, -0.1156000, -0.2004540, 0.0903189, 0.1912550, 0.0491491, 0.2571260, 0.3284450, 0.0962949, -0.0437188, -0.1510300, 0.1461060, 0.1488620, 0.1929070, -0.1042680, -0.2973560, -0.2182430, -0.2812070, -0.0728197, -0.0046743, 0.1678340, 0.0938065, 0.1359640, 0.0409524, 0.0088634, -0.0002811, -0.0002272, 0.0168263, -0.0481147, -0.0589850, -0.1304870, -0.0214897, 0.0060140, 0.1166660, 0.2221610, 0.1955210, 0.0058101, -0.0728106, -0.0365949, 0.0654353, 0.0154690, -0.1240430, -0.3755790, -0.2060420, -0.1893780, -0.0951864, -0.0197494, 0.0993535, 0.1924490, 0.1010300, 0.1212650, 0.0185542, -0.0012856, 0.0022427, -0.0000433, -0.0066190, -0.0884590, -0.0019353, -0.1697070, -0.1624990, -0.0382805, -0.1177190, -0.0799640, 0.0067605, -0.1271760, -0.0393191, -0.1066700, -0.1460010, -0.3670780, -0.3283020, -0.2256050, -0.0398612, 0.1092840, 0.1212040, 0.1096670, 0.2410570, 0.2942370, 0.1225190, 0.0523609, 0.0108217, -0.0037252, 0.0000050, 0.0010329, -0.0049838, -0.1398240, -0.0797227, -0.1305790, -0.1765970, -0.1456100, -0.2707700, -0.1687260, 0.0236955, -0.1957440, -0.4868080, -0.4743820, -0.3936950, -0.2936000, -0.1717280, -0.0149555, -0.0005323, 0.1796930, 0.1371870, 0.2246310, 0.2538440, 0.1573040, 0.0496954, 0.0053983, 0.0040298, -0.0010478, 0.0004252, -0.0013939, 0.0026760, -0.0327365, -0.0227495, -0.0597667, 0.0821124, 0.0655047, -0.1053820, -0.1615780, -0.0758410, -0.2496040, -0.3217350, -0.4367360, -0.3607580, -0.1469440, -0.0750497, -0.1259260, -0.0223139, 0.0776725, 0.2613070, 0.3211880, 0.2044600, 0.1067090, 0.0456000, 0.0002487, 0.0002875, -0.0002169, 0.0005825, 0.0007909, 0.0493618, 0.0707886, 0.1912230, 0.1160770, 0.1587660, 0.0579498, 0.0107181, -0.0713915, -0.1020200, -0.0962103, -0.2899730, -0.1079780, -0.0747077, 0.0506208, 0.0850019, 0.0314498, -0.0704854, 0.2397490, 0.2236510, 0.2244780, 0.1898420, 0.0905409, 0.0263871, 0.0036554, -0.0194516, 0.0001511, 0.0003404, -0.0004635, 0.0520194, 0.1014770, 0.2017170, 0.2239600, 0.1889300, 0.2348680, 0.1536000, -0.0994883, -0.0179262, -0.0108067, 0.0213823, -0.0539598, -0.0522388, -0.0014524, 0.0989353, 0.0749569, 0.1538530, 0.2863160, 0.2357910, 0.1364960, 0.0828163, 0.0542815, 0.0285347, 0.0040660, -0.0037147, 0.0002256, 0.0004514, 0.0001716, -0.0085042, -0.0045878, 0.0417022, -0.0138554, 0.0670866, 0.1125350, 0.1515420, -0.0701671, -0.2337420, -0.1209490, -0.0670727, 0.1841300, 0.0949674, 0.2263050, 0.1354320, 0.1666860, 0.2151100, 0.1955140, 0.1165090, 0.0754934, 0.0600333, 0.0265553, 0.0048540, -0.0030139, -0.0025460, 0.0006532, -0.0004109, -0.0001094, 0.0000669, -0.0065012, -0.0176416, -0.0553495, 0.1039430, 0.1035080, 0.0517516, 0.1037250, 0.2298580, 0.2959650, 0.1828400, 0.1703620, 0.1151630, 0.1033880, 0.0666950, -0.0532318, 0.0126143, 0.0426785, 0.0619043, 0.0696181, 0.0315805, 0.0087149, 0.0006235, 0.0007142, -0.0001618, -0.0001011, 0.0002967, -0.0000327, -0.0003703, -0.0003844, -0.0052188, -0.0116946, 0.0484617, 0.0811217, 0.0830458, 0.0706524, 0.2775120, 0.2925560, 0.2618430, 0.2221950, 0.2220370, 0.1676970, 0.0586351, 0.0320526, 0.0283501, 0.0315857, 0.0230521, 0.0050742, 0.0004656, -0.0017084, -0.0009543, -0.0002966, 0.0000024, 0.0001646, -0.0001271, -0.0003610, 0.0001369, 0.0000855, 0.0005403, -0.0023422, 0.0225354, 0.0494124, 0.0618320, 0.0800138, 0.0812283, 0.0542974, 0.0485649, 0.0496095, 0.0330888, -0.0147419, -0.0311997, -0.0117983, 0.0085964, 0.0032590, 0.0036591, 0.0020955, 0.0015206, 0.0001389, -0.0001317, -0.0001846, 0.0000400, 0.0000042, -0.0002886, 0.0002465, 0.0003870, 0.0002595, 0.0003759, 0.0001243, 0.0000533, 0.0030340, 0.0032711, 0.0035611, 0.0068940, 0.0043018, 0.0036371, 0.0073595, 0.0064550, 0.0017124, 0.0062582, 0.0037771, 0.0030239, 0.0013538, 0.0003321, -0.0000536, 0.0010449, -0.0000042, -0.0001647, -0.0001166, -0.0001889, -0.0001038, -0.0000200, 0.0001379, 0.0004640, -0.0001158, -0.0007763, 0.0002835, -0.0003408, 0.0000400, 0.0000659, -0.0004205, -0.0004031, -0.0004197, 0.0011812, 0.0040291, 0.0001467, -0.0004091, 0.0000887, -0.0005639, -0.0002107, -0.0004664, -0.0006183, 0.0000107, -0.0000857, 0.0004035, 0.0000534, -0.0001628, -0.0001707, 0.0001811, 0.0006446, -0.0007829, -0.0000100, -0.0003189, -0.0001820, -0.0001393, 0.0123128, 0.0217222, 0.0269396, 0.0141298, 0.0306823, 0.0267616, 0.0380749, 0.0522883, 0.0316933, 0.0238961, 0.0182311, 0.0192408, 0.0270676, 0.0270004, 0.0334304, 0.0289718, 0.0146817, 0.0065773, 0.0005268, 0.0000291, -0.0001831, 0.0002159, 0.0007325, 0.0001083, 0.0005557, 0.0000249, 0.0018251, 0.0011352, 0.0165522, 0.0457060, 0.0469968, -0.0077859, -0.0067627, 0.0480638, 0.0645408, 0.0411421, 0.0645891, 0.0415407, 0.0678978, 0.1115470, 0.1392340, 0.1456480, 0.0986603, 0.0567067, 0.0232349, 0.0197081, 0.0015771, -0.0014120, 0.0000558, -0.0005922, 0.0002837, -0.0004298, -0.0060174, 0.0035717, 0.0252948, -0.0047168, 0.0134785, -0.0046520, -0.0304744, -0.0555244, -0.1134990, -0.1447720, -0.1448260, -0.0070760, 0.0004793, 0.0238549, -0.0268490, 0.1461970, 0.2669060, 0.3304810, 0.2256730, 0.2228650, 0.0739837, 0.0271765, 0.0366876, 0.0079154, 0.0179896, -0.0004810, 0.0002232, 0.0000196, -0.0207637, -0.0037890, -0.0015479, -0.0976886, -0.1328620, -0.1085030, -0.1721740, -0.1648720, -0.1322090, 0.0006211, -0.1491060, -0.0438832, 0.0656866, 0.0041501, -0.0053106, 0.0616037, 0.0124056, 0.1081810, 0.1628920, 0.1825790, 0.0917998, 0.2820010, 0.1764230, 0.0775820, 0.0095682, 0.0009075, 0.0000444, -0.0002575, -0.0027723, 0.0014475, -0.0856147, -0.0748747, -0.0779972, -0.1465070, 0.0212142, -0.0261164, -0.0375298, -0.0164195, 0.0027071, -0.0586514, -0.1058490, -0.1889400, -0.0334934, -0.0031518, 0.0061777, -0.0972037, 0.2232090, 0.1258260, 0.2723540, 0.3122180, 0.1292990, 0.0301786, 0.0043846, 0.0041519, 0.0000936, 0.0001125, 0.0173568, -0.0533693, -0.1658050, -0.0421792, -0.1890970, -0.0850146, 0.0453209, -0.0414976, 0.0137934, -0.0844122, -0.0129463, -0.0964799, 0.1251290, 0.1683720, -0.0106795, 0.2593620, 0.3581690, 0.1118020, 0.2645280, 0.1219360, 0.2368300, 0.1509550, 0.1596010, 0.0632519, 0.0233033, 0.0096926, -0.0003462, -0.0056153, 0.0073767, -0.1209710, -0.2182370, -0.0805273, -0.1766660, 0.0408467, 0.1120810, 0.1466760, 0.2281680, 0.0708960, 0.1329670, 0.1345040, 0.3052050, 0.2937160, 0.4064040, 0.5005090, 0.4948980, 0.3771980, 0.4250680, 0.3241000, 0.2109690, 0.0943515, 0.0995467, 0.0707787, 0.0175275, 0.0066916, -0.0012008, -0.0003158, -0.0019299, -0.0733537, -0.2035360, -0.1575930, -0.0563152, -0.0568919, 0.0538568, -0.0323117, -0.2215240, 0.0775731, 0.0834689, 0.0401062, -0.0377032, 0.1508430, 0.1621020, 0.1286290, 0.2884280, 0.3313630, 0.2262860, 0.0173874, 0.0017799, -0.0261489, 0.0097252, -0.0140583, 0.0010577, 0.0091194, 0.0003182, 0.0000318, -0.0052172, -0.0492820, -0.1454180, -0.1835860, -0.1675390, -0.2051690, -0.0642887, -0.0790917, -0.1365930, -0.0953384, -0.2496710, -0.3482470, -0.3074770, -0.4040870, -0.6640480, -0.7842220, -0.7408610, -0.6045830, -0.6197880, -0.4056230, -0.5076700, -0.6002900, -0.2555500, -0.1555970, -0.0277318, 0.0001468, 0.0000785, 0.0001520, -0.0023469, -0.0478802, -0.0385214, -0.1855020, -0.0936332, -0.1533190, -0.0104348, 0.1089640, -0.2224890, -0.1307780, -0.2349100, -0.1587360, -0.5414890, -0.4125030, -0.7203540, -1.2438900, -1.2663200, -1.2777100, -1.0875300, -0.8412800, -0.7506560, -0.7112560, -0.3244330, -0.1553320, -0.0180357, -0.0005576, -0.0000243, -0.0006874, -0.0015877, -0.0391562, -0.0104802, -0.0445466, 0.1274630, -0.0010127, -0.1334400, -0.1613040, -0.0024472, -0.1106320, -0.1881210, -0.0553723, -0.0926368, 0.0119347, -0.0532961, -0.2866510, -0.3058220, -0.5814010, -0.6358860, -0.5028050, -0.5554680, -0.5172660, -0.3606660, -0.1418500, -0.0262651, 0.0028746, 0.0003519, -0.0001228, -0.0006801, -0.0087045, -0.0059371, -0.0659825, 0.0363316, 0.0058294, 0.1008670, 0.0732451, 0.0187818, 0.0450727, -0.0715791, -0.1399340, -0.1628900, 0.1070670, 0.0535646, 0.0313040, 0.1731240, -0.0060666, 0.0846939, -0.0050168, -0.1719430, -0.2017840, -0.1991440, -0.1526960, -0.0125129, 0.0031315, -0.0003537, 0.0003801, 0.0015445, -0.0429742, -0.0089867, -0.1139970, 0.0953501, 0.1102660, -0.1878240, 0.0212390, 0.1049770, -0.0447456, -0.0988414, 0.0137775, 0.0770205, 0.1218180, -0.0200981, 0.0056014, 0.1801370, 0.1334630, 0.0923597, 0.0201591, -0.0254662, -0.1048000, -0.1380200, -0.1229690, -0.0392560, -0.0044243, 0.0002841, -0.0010856, 0.0003131, -0.0545762, -0.0354049, -0.1405800, 0.0180920, 0.0990526, -0.0791581, -0.0757517, 0.0356220, 0.0830898, -0.0033241, -0.0965880, -0.0024894, 0.0618922, 0.1602090, -0.1186130, 0.3126890, 0.0491296, 0.2246680, -0.0460311, 0.0014404, -0.0388652, -0.0996685, -0.0929985, -0.0427441, -0.0002211, 0.0003108, -0.0034777, -0.0059638, -0.0687337, -0.1547820, 0.0451566, 0.0853153, 0.0378651, -0.0012019, -0.0870374, 0.1109310, -0.0936751, 0.1015800, 0.0106206, -0.0337090, -0.0245230, 0.1430610, 0.0561410, 0.2421690, 0.0318113, 0.1031340, -0.0794440, -0.1873170, 0.0140849, 0.0784730, -0.0294045, -0.0821843, -0.0158755, -0.0001653, -0.0024702, -0.0148544, -0.0542907, -0.1703460, -0.0542372, -0.0543792, -0.0495060, 0.0316904, -0.1495790, -0.0354166, 0.0040794, 0.0697249, 0.1618260, 0.0856532, 0.1655650, 0.2686920, 0.1972260, 0.0509941, -0.1048810, -0.0855826, -0.1485590, -0.0298434, -0.1411880, 0.0744089, -0.0433316, -0.1014520, -0.0389021, 0.0004547, -0.0003309, -0.0304904, -0.0234622, -0.1523700, -0.0903610, 0.0509740, -0.0614964, 0.0460086, -0.1054150, 0.0749102, -0.0437724, 0.1249340, -0.1308190, -0.0068384, 0.1979800, -0.0110177, -0.0029567, 0.0455868, -0.0202617, 0.1573650, 0.0766482, 0.1437640, 0.0292615, 0.1949110, -0.0123435, -0.0151669, -0.0135241, 0.0004385, -0.0002116, -0.0235664, -0.0475273, -0.0512729, 0.0517451, -0.0836578, 0.0816072, -0.0304437, 0.0664483, 0.1468350, -0.2075640, 0.2021770, -0.0272291, 0.2825380, 0.1784410, 0.0041848, -0.0204574, 0.0894626, 0.0268200, 0.1080950, 0.0064470, 0.0068716, -0.0533622, 0.1227180, 0.0308293, 0.0146250, -0.0057745, -0.0000635, -0.0000907, 0.0373734, -0.0414775, 0.0037813, 0.0646805, 0.0000650, -0.0714841, 0.0994451, 0.0651626, 0.0710772, 0.1195770, 0.2013650, 0.1273610, 0.1892320, 0.0474052, -0.0272691, -0.0656026, 0.0579802, 0.0722656, -0.0286489, -0.0224677, 0.0182956, 0.0175491, 0.1299550, 0.0369587, -0.0221492, -0.0020570, 0.0000457, -0.0008766, 0.0376418, -0.0199062, 0.1440480, 0.1620970, -0.0354098, -0.2501690, 0.0479941, -0.0713049, 0.0096818, 0.0621400, -0.0952886, 0.0714670, 0.1093870, 0.1234630, -0.0262371, -0.1122270, 0.0992751, 0.1126920, -0.1099490, 0.0416437, 0.0649314, 0.0797085, 0.1053680, 0.0947144, -0.0079279, 0.0008389, 0.0001381, -0.0007265, -0.0101887, -0.0176380, 0.1714410, 0.1449360, 0.0104781, -0.0399660, -0.2173000, -0.1948910, 0.0826821, -0.0359844, 0.1263680, 0.1985470, 0.2162140, 0.0569804, 0.1630660, 0.0402271, 0.0012067, -0.0542719, 0.1363180, 0.1934980, 0.1131240, 0.0445369, 0.1454140, 0.1009690, 0.0000238, -0.0000471, -0.0003418, 0.0004239, -0.0076765, -0.0006829, 0.1030630, -0.0038542, -0.0428497, -0.1489070, -0.0802112, -0.0032941, 0.0735562, 0.0217971, 0.1986560, -0.0311494, 0.0535668, 0.0796800, 0.0361291, 0.0969398, -0.0198956, -0.0746146, 0.0522072, -0.0470636, -0.0364203, 0.0086829, 0.0510781, 0.0488471, 0.0099017, 0.0000502, -0.0000835, -0.0000543, -0.0159532, -0.0417598, 0.0462743, 0.0508341, 0.0466694, -0.1519170, -0.1294800, 0.0106297, 0.1180200, -0.2471290, -0.1326900, -0.1109390, 0.0382395, 0.0075505, 0.0775622, -0.1001560, -0.1638930, -0.0162933, 0.0623109, -0.0258495, -0.0408405, -0.0667498, 0.0062062, 0.0265114, 0.0042074, 0.0001644, -0.0002813, -0.0002919, -0.0125523, -0.0534627, -0.0719890, -0.0246658, -0.0588214, -0.1664810, -0.2467770, -0.1066920, -0.0074649, -0.1278670, 0.0455534, 0.1308240, 0.0859109, 0.1708600, -0.1756440, -0.1715080, -0.0144668, -0.0721505, -0.0189418, -0.0603632, -0.0616704, -0.0602192, -0.0186607, -0.0082027, -0.0002576, 0.0004618, 0.0000877, -0.0000122, -0.0017666, 0.0007496, -0.0205406, -0.0477971, -0.0495883, -0.0602230, -0.0902777, -0.0061475, -0.1305790, -0.0053072, 0.3062530, 0.1863160, 0.1295390, 0.1942360, 0.0618033, 0.0043927, 0.0596160, 0.0786943, -0.0170728, 0.0188550, 0.0398714, 0.0114616, 0.0060522, -0.0006706, -0.0001313, 0.0001352, 0.0002115, -0.0000363, -0.0004669, 0.0006700, -0.0007139, 0.0000356, 0.0048287, 0.0115697, 0.0095192, 0.0143067, 0.0114701, 0.0196408, 0.0027073, 0.0857469, 0.1101490, 0.1410250, 0.0955007, 0.0598965, 0.0219925, 0.0335810, 0.0322652, 0.0284649, 0.0118969, 0.0008078, 0.0001554, -0.0001204, -0.0002336, -0.0000206, 0.0004662, 0.0004580, 0.0003313, 0.0004379, -0.0001368, -0.0000587, -0.0004853, 0.0002253, -0.0001375, 0.0004696, 0.0003577, 0.0002889, 0.0002806, 0.0007110, 0.0006112, -0.0007242, 0.0003810, -0.0004739, 0.0009922, 0.0006149, -0.0001858, -0.0063396, -0.0036363, 0.0004770, 0.0003015, 0.0003020, -0.0000513, 0.0005530, -0.0007597, 0.0000937, -0.0005398, 0.0002306, -0.0000418, 0.0003503, -0.0000593, 0.0000573, -0.0004927, 0.0004746, 0.0006073, 0.0002274, 0.0001784, 0.0002621, -0.0005226, 0.0005796, -0.0001486, 0.0005549, 0.0006013, 0.0011091, 0.0001937, 0.0003766, 0.0006426, 0.0000603, 0.0005388, 0.0004715, -0.0008365, -0.0002315, 0.0001780, 0.0002895, 0.0000003, -0.0004184, 0.0004410, 0.0005016, -0.0004128, -0.0004363, -0.0006913, -0.0003117, -0.0029313, -0.0015001, -0.0003554, -0.0007964, 0.0015112, 0.0012101, -0.0031935, -0.0012082, 0.0000027, -0.0010410, -0.0014484, -0.0003522, -0.0002161, 0.0001813, 0.0000805, 0.0000212, 0.0000626, 0.0000835, 0.0001877, -0.0000472, -0.0004984, -0.0004761, 0.0005211, -0.0005729, 0.0001964, -0.0010017, -0.0015806, 0.0096048, 0.0021160, 0.0017592, 0.0020053, 0.0203874, 0.0328393, 0.0324555, 0.0279146, 0.0191888, -0.0050698, 0.0042680, 0.0197000, 0.0150289, 0.0042387, 0.0021858, 0.0014966, 0.0001419, 0.0003268, -0.0005434, -0.0005104, 0.0002350, 0.0002248, -0.0004804, -0.0025851, 0.0093883, 0.0101269, 0.0248252, 0.0160594, -0.0303937, -0.0488293, -0.0217809, -0.0392443, 0.0384491, 0.1087730, 0.0958836, 0.1147310, 0.0747000, 0.0836074, 0.0516111, 0.0662692, 0.0097155, 0.0127863, 0.0577605, 0.0476471, -0.0440623, -0.0129649, 0.0005314, 0.0000853, -0.0001601, -0.0001062, 0.0002746, 0.0002102, 0.0315109, 0.0526253, 0.0663700, 0.0539289, 0.0001373, 0.0193824, -0.0005494, 0.0338317, 0.0573170, -0.0323370, 0.0144985, 0.0916082, 0.0266290, 0.1292570, 0.2023280, 0.1611210, 0.1397350, 0.2143190, 0.0641702, -0.0072241, -0.0362807, -0.0036683, 0.0005589, 0.0003388, 0.0001637, 0.0000927, 0.0010966, -0.0362186, -0.0233362, 0.0069388, 0.0463354, 0.0440524, 0.1145670, 0.2960820, 0.1751170, 0.2769520, 0.1886630, 0.1057310, 0.2133270, 0.2864120, 0.3625180, 0.4169130, 0.4176070, 0.3265180, 0.2028700, 0.1793320, 0.1444490, 0.0442578, -0.0185783, -0.0088754, 0.0012372, 0.0001474, -0.0002543, -0.0112587, -0.0209754, -0.1034290, -0.0946468, -0.0737397, -0.0020258, 0.0048621, 0.0912160, 0.1483190, 0.0286653, 0.1639800, 0.1603760, 0.2611420, 0.4309560, 0.5071900, 0.4086830, 0.4874050, 0.4489870, 0.3416080, 0.1450760, 0.0323359, 0.0671938, -0.0646069, -0.0329036, -0.0408325, 0.0001511, -0.0007508, -0.0023456, -0.0126011, -0.0327436, -0.0356109, -0.0270674, -0.0248479, -0.0500140, -0.0712540, -0.0876273, -0.0721276, 0.1345470, -0.0648063, 0.0180741, 0.0533883, -0.0226850, -0.0373503, -0.1646210, -0.0667458, -0.0179598, -0.2595700, -0.0999397, -0.1057040, -0.0511331, -0.0280351, 0.0058439, -0.0423572, -0.0008964, 0.0013243, -0.0152025, -0.0121286, -0.0124923, 0.0479390, -0.0217633, -0.0872897, -0.0576876, -0.2618000, -0.1915000, -0.0749227, -0.1612590, -0.0871138, -0.1016420, -0.1778410, -0.4408470, -0.4751350, -0.4728320, -0.4639790, -0.2147890, -0.3387000, -0.2000830, -0.2260230, -0.2122820, -0.1736320, 0.0045919, -0.0057082, -0.0023097, -0.0004625, -0.0162211, -0.0214573, -0.0081274, 0.0404544, 0.0247448, -0.0444287, 0.0288453, -0.1509760, -0.1480400, -0.2095980, -0.2779330, -0.3339310, -0.1752220, -0.3652240, -0.3233990, -0.4316520, -0.5917450, -0.5807040, -0.4146290, -0.1814020, -0.1813360, -0.2013580, -0.1133030, -0.0954103, -0.0487507, -0.0459623, -0.0378885, -0.0003031, -0.0138921, -0.0248930, 0.0175646, 0.0112403, -0.0408951, -0.0478109, 0.0800386, -0.1010440, -0.2718610, -0.2490690, -0.2199030, 0.0159326, -0.3361430, -0.2614260, -0.1847590, -0.4235240, -0.1266260, -0.2841670, -0.1556080, -0.0554571, -0.0287408, -0.0524444, -0.0733950, -0.1245070, -0.0890013, -0.0518269, -0.0104751, -0.0005251, -0.0080534, -0.0473367, 0.0031441, -0.0057409, 0.0052464, -0.0110426, -0.0476394, -0.1488890, -0.0502132, 0.0283749, -0.2535450, -0.1981900, -0.1917890, -0.0328021, -0.1711080, -0.0156208, 0.3206500, 0.1221680, 0.1505060, 0.2216800, 0.1065810, -0.1374140, -0.1566130, -0.1409680, -0.0803533, -0.0413866, -0.0033331, 0.0000613, -0.0041515, -0.0395408, -0.0241090, -0.0837580, 0.0621945, 0.0311218, -0.1505020, -0.0595908, -0.0693200, 0.1144470, -0.0336419, 0.0260893, -0.0677837, -0.0006350, -0.1047450, 0.3905750, 0.4885550, 0.2048090, 0.1431010, 0.1715640, 0.1605370, -0.1054680, -0.1745250, 0.0140340, -0.0613186, -0.0644993, -0.0041946, -0.0000276, -0.0025663, -0.0236777, -0.0068858, -0.0251773, -0.0674416, 0.0297321, 0.0575269, 0.0783257, 0.0031474, 0.0636001, 0.0164201, -0.0040548, 0.0627596, -0.0498493, 0.0198742, 0.2393640, 0.4547250, 0.3305570, 0.1167290, 0.0747371, -0.0778583, -0.0487223, -0.0139444, -0.0235335, -0.0380528, -0.0264845, 0.0037928, -0.0008092, -0.0017010, -0.0155139, 0.0011916, 0.0470820, 0.0100997, 0.1067300, 0.1064440, 0.0703848, 0.0153041, -0.0966830, -0.0140595, 0.0121600, 0.0709167, -0.0150614, 0.0619208, 0.0673661, 0.0759359, -0.0354612, 0.1050470, -0.0430948, -0.0461825, -0.0054867, 0.0045169, -0.0205511, 0.0283086, -0.0037008, -0.0000195, -0.0002620, -0.0001397, -0.0015936, 0.0482969, 0.0717633, -0.0155014, -0.0129041, 0.0293649, 0.1023510, -0.0051296, -0.0244350, -0.0531172, 0.0829277, 0.2666320, 0.0689207, 0.1592840, 0.2484650, -0.0052500, -0.1629200, -0.0230263, 0.0401332, -0.0881685, 0.0513290, -0.0850953, -0.0161944, 0.1059450, 0.0601279, 0.0055740, 0.0004123, 0.0008711, -0.0024628, 0.0797988, 0.1036920, -0.0466085, -0.0713808, -0.0157714, -0.0731016, 0.0192986, -0.1345660, -0.0461891, 0.2012840, 0.3006440, 0.2623850, 0.3112170, 0.0766365, -0.0270976, -0.0089754, 0.0446658, 0.1261930, 0.0342170, 0.0383912, 0.0116757, 0.0769980, 0.1299230, 0.0417079, 0.0104687, 0.0002579, 0.0001596, 0.0022961, 0.0292524, 0.1298720, -0.0333989, -0.0860638, -0.0253424, -0.1402610, -0.1065930, -0.1201560, 0.1018960, 0.4683840, 0.3143800, 0.0301964, -0.1416850, -0.0239020, -0.1192180, 0.1022920, 0.0301488, -0.0381898, 0.1035580, 0.0165928, 0.0122877, -0.0395252, 0.0645839, 0.0013706, 0.0006089, -0.0013385, 0.0005447, 0.0031259, 0.0538157, 0.1613720, 0.0695027, -0.0057133, -0.0832004, -0.1176180, -0.1181080, 0.0439018, 0.1442750, 0.0651370, 0.0272638, -0.1066630, 0.1702640, 0.0902290, -0.0623103, 0.1263200, 0.0334039, -0.0176025, 0.1934390, 0.0503543, 0.0671958, 0.0234795, 0.0303148, -0.0088891, 0.0005884, -0.0001130, -0.0066132, 0.0034155, 0.0969005, 0.0856383, 0.0799414, -0.0032903, 0.0726823, -0.0466736, 0.0565293, 0.0573353, 0.0834123, -0.1081190, 0.0188683, -0.0132575, 0.0711117, 0.1853600, -0.0947785, 0.1175240, -0.0360122, 0.0770994, 0.1728060, 0.1676070, 0.0694989, -0.0083333, -0.0076669, 0.0133872, -0.0002015, -0.0001872, -0.0014813, 0.0095384, 0.1177410, 0.1685860, 0.0769596, 0.0592102, 0.1996120, -0.0330852, -0.0392485, -0.0518114, 0.0041582, -0.0056521, 0.0167426, 0.0266499, 0.1622310, 0.2741730, 0.0164564, 0.1715460, 0.0865104, 0.0822274, 0.1479370, 0.1395480, 0.0349381, -0.0817918, -0.0677365, 0.0055737, -0.0000897, -0.0005890, 0.0000228, 0.0121607, 0.0897133, 0.1209340, 0.0833044, 0.1244390, 0.1501040, 0.0488594, -0.1792680, -0.0218213, -0.0416239, -0.0026542, 0.0099704, 0.0588131, 0.1258150, 0.0893574, -0.0359606, 0.0711532, 0.0462607, 0.0878900, 0.1051610, 0.1153040, 0.0250059, -0.0835261, -0.0797198, 0.0007002, -0.0002651, 0.0002081, -0.0006427, 0.0094360, 0.0132975, 0.0369232, 0.0685503, 0.1361890, 0.0773817, 0.0917305, -0.0133027, 0.0582825, 0.1822860, -0.0478243, 0.0830925, 0.0235057, -0.0733840, -0.1207150, -0.0320465, 0.0991266, 0.1705920, 0.0220247, 0.0981070, 0.0684466, 0.0068413, -0.0770107, -0.0517038, 0.0006114, -0.0003340, 0.0004050, -0.0001292, 0.0155821, 0.0075753, -0.0206598, -0.0165959, 0.0084879, -0.0023115, 0.0653298, 0.1531590, 0.0702733, 0.0719944, -0.0114578, 0.0306497, 0.0450522, 0.0138738, -0.1896270, 0.0912851, 0.1751830, 0.1143480, 0.0325066, 0.0983698, 0.0361818, -0.0285116, -0.0499377, -0.0153976, 0.0029293, 0.0000789, -0.0005293, -0.0002534, 0.0110530, 0.0097574, -0.0167884, -0.0688831, 0.0624332, 0.0884952, 0.1037590, 0.1888860, -0.0531709, -0.0090652, -0.0405743, 0.0851651, 0.0732457, -0.0825626, -0.0757110, 0.0192334, 0.1392900, 0.0136747, -0.0013196, 0.0355951, 0.0072519, -0.0257942, -0.0112459, 0.0133623, 0.0002097, -0.0001759, -0.0000049, 0.0007128, 0.0016102, -0.0060019, -0.0326841, -0.0571665, -0.0081303, -0.0162245, 0.0504199, 0.1026250, 0.0664302, -0.0825291, -0.1122110, 0.0247675, 0.0574792, 0.0051872, -0.1391220, -0.1929600, -0.1088250, -0.1675730, -0.0475488, -0.0609562, -0.0549994, -0.0378712, -0.0239606, 0.0002276, 0.0003852, 0.0002393, -0.0004259, -0.0003670, 0.0007246, 0.0002286, 0.0002758, -0.0016388, -0.0195002, -0.0408672, -0.0688402, -0.1046890, -0.0505841, -0.0640761, -0.0838037, -0.1886850, -0.1208990, -0.0559288, -0.0571235, -0.0287599, -0.0707376, -0.1239090, -0.0746232, -0.0285132, -0.0208128, -0.0028694, -0.0013048, 0.0004449, 0.0000994, 0.0001023, -0.0001843, 0.0002444, 0.0001778, -0.0001797, -0.0003843, 0.0002818, -0.0006411, -0.0052877, -0.0047264, -0.0013380, -0.0160544, -0.0041603, -0.0064618, -0.0066568, -0.0079230, 0.0157881, -0.0025309, -0.0124857, -0.0305713, -0.0193469, -0.0101411, -0.0012214, -0.0092774, -0.0034052, -0.0001576, 0.0002123, 0.0004124, -0.0000698, -0.0004331, 0.0004365, 0.0001359, 0.0003083, -0.0001677, 0.0000404, 0.0003204, 0.0001894, -0.0000493, -0.0000239, -0.0003497, -0.0005566, 0.0000752, -0.0000794, -0.0004955, 0.0003053, 0.0001128, -0.0001949, -0.0005811, -0.0002147, 0.0000222, -0.0003351, 0.0000828, -0.0000134, -0.0000361, -0.0001221, 0.0004129, -0.0002344, -0.0001423, -0.0004148, -0.0003045, -0.0002221, -0.0003707, -0.0000309, -0.0000907, -0.0007147, -0.0022777, -0.0034542, -0.0020518, -0.0001610, -0.0011978, -0.0033178, 0.0192435, 0.0389326, -0.0266568, -0.0087487, -0.0013427, -0.0022375, -0.0008833, 0.0027745, -0.0002665, 0.0002743, 0.0000850, 0.0000227, -0.0003733, 0.0000041, 0.0004626, 0.0000097, 0.0000278, -0.0002110, 0.0002000, -0.0001542, 0.0006357, -0.0004599, -0.0047561, -0.0116354, -0.0094375, -0.0089167, -0.0300407, -0.0731649, -0.0912920, -0.0936369, -0.0880888, -0.0476896, -0.0141506, -0.0304741, -0.0371283, -0.0175812, -0.0086086, -0.0079502, -0.0047701, -0.0017072, -0.0002971, -0.0001004, 0.0006392, 0.0000340, 0.0011866, 0.0009347, 0.0071072, 0.0017537, 0.0012056, 0.0120674, -0.0109336, -0.0186307, -0.0068332, -0.0472945, -0.1750540, -0.4185760, -0.4796100, -0.3168010, -0.2407370, 0.0122799, -0.0057477, 0.0941405, 0.1112940, 0.0353995, 0.0387841, -0.0278292, -0.0297052, -0.0034335, -0.0087726, -0.0001551, 0.0003403, -0.0002371, 0.0052710, 0.0010537, -0.0027248, 0.0022615, 0.0022663, 0.0055693, 0.0001199, -0.0024535, -0.0653383, -0.1959470, -0.3591250, -0.5437830, -0.3172900, -0.0618424, 0.0345264, 0.0789420, -0.0668211, 0.0467006, 0.0630357, -0.0919966, -0.0745194, -0.0100004, -0.1106720, -0.0594336, -0.0202473, -0.0064257, -0.0000275, 0.0001856, 0.0004546, 0.0096315, -0.0014666, 0.0143369, 0.0346312, 0.0571831, 0.0189809, -0.0330661, -0.2074070, -0.5798520, -0.7920150, -0.5747000, 0.0107812, 0.0486482, 0.0811018, 0.0690579, -0.2052190, -0.2111320, -0.0822038, -0.0260707, 0.0279259, 0.0260272, 0.0039965, -0.0883373, -0.0241506, -0.0045557, 0.0002382, -0.0000365, -0.0112146, -0.0205057, -0.0355987, 0.0630712, 0.1422940, 0.0984891, 0.0755135, 0.0543485, -0.1986740, -0.6679040, -0.8644730, -0.6911160, -0.0210423, 0.0965508, 0.0693700, -0.0335836, -0.1312960, -0.1640320, 0.0847347, -0.0624351, 0.0334174, 0.1437340, -0.0121311, -0.0717451, 0.0144301, -0.0001705, -0.0003703, -0.0003238, -0.0087365, -0.0277770, 0.0516896, 0.1925390, 0.1090680, 0.0808659, 0.0589994, 0.1373620, -0.1441910, -0.6341370, -0.8168330, -0.4235310, 0.2830440, 0.3068210, 0.1506520, 0.0717027, -0.2435770, -0.0409845, 0.0253395, 0.0830975, 0.1368970, 0.0383634, -0.1763520, -0.1378570, 0.0175589, -0.0053741, 0.0015473, -0.0048383, -0.0044686, -0.0108286, 0.0734292, 0.1622660, 0.0622636, -0.0286439, 0.0501852, 0.1386610, -0.1493150, -0.6548040, -0.8934020, -0.2870650, 0.1758100, 0.4178580, 0.0872940, 0.2697640, -0.1373250, 0.0120399, -0.0316120, -0.0624292, -0.0444730, -0.1050040, -0.0521754, 0.0037712, -0.0057608, -0.0000138, -0.0006254, -0.0079760, -0.0070369, -0.0209199, 0.0684322, 0.1088670, 0.0078288, 0.0197209, 0.1411500, 0.1015850, -0.0970885, -0.6196470, -0.8551810, -0.2424570, -0.0085460, 0.3897980, 0.4028350, 0.3247370, 0.1335190, 0.0962236, -0.1462640, -0.0564155, -0.1737610, -0.0606000, 0.0759777, 0.0044629, 0.0431127, 0.0021161, 0.0000131, -0.0056534, -0.0078742, -0.0266328, 0.0450161, 0.0203129, -0.0365937, 0.1158770, 0.1596140, 0.0233970, -0.1488780, -0.6214660, -0.5077730, -0.2079120, 0.0759745, 0.5507610, 0.3580440, 0.3504140, 0.1519760, 0.0464720, -0.0875078, -0.0233933, -0.1075820, 0.0356131, 0.1415710, 0.1606930, 0.0312879, 0.0003175, 0.0000218, -0.0042283, -0.0222674, -0.0240947, -0.0117766, -0.0225409, -0.0314276, -0.0088111, 0.0584804, -0.0309186, -0.1992460, -0.4234070, -0.2030340, 0.0639187, -0.0419047, 0.2766700, 0.3040650, 0.2123340, 0.0284765, -0.2138510, -0.0821513, 0.0629524, -0.0651524, 0.0239104, 0.0878488, 0.0787457, -0.0278258, -0.0013617, -0.0003815, -0.0021666, -0.0224886, -0.0222260, -0.0568085, -0.0948470, 0.0380774, -0.0623290, -0.0146611, 0.0420734, -0.0615897, -0.1708200, 0.1435830, 0.0236844, -0.0303455, 0.0817443, 0.2270020, -0.0335436, -0.0633291, -0.2491460, -0.0410510, 0.0946715, 0.0175336, -0.0895000, -0.0427410, 0.0205439, -0.0166276, -0.0035982, 0.0004439, -0.0030765, -0.0188756, -0.0199386, -0.0919049, -0.1036060, 0.0611078, -0.0208795, -0.0721434, 0.0123633, -0.0295152, 0.0269641, 0.1641140, 0.0407347, -0.0094860, -0.1846660, 0.0537664, 0.0786698, -0.1068420, -0.1896870, -0.1287870, -0.0318258, -0.1096480, -0.1070810, -0.0859471, -0.0295153, -0.0195458, -0.0014122, -0.0002598, -0.0023954, -0.0083089, -0.0118335, -0.0425338, -0.0823493, -0.0331553, 0.0480482, 0.1430860, 0.1174670, -0.0048767, 0.1489290, 0.0765046, -0.0772534, 0.0163746, 0.0360747, 0.2471100, 0.0950359, -0.1102800, 0.0034273, -0.1304170, -0.0023857, -0.0391950, -0.1118610, -0.0119817, -0.0072148, -0.0006884, 0.0000081, -0.0001218, -0.0006927, -0.0004787, -0.0248030, 0.0165492, -0.0889524, -0.0599434, 0.2627730, 0.1655230, 0.1304250, -0.0840989, 0.0074014, -0.0109808, 0.0194535, -0.1362710, -0.1080110, 0.0184972, -0.0582773, -0.0533403, -0.0639651, -0.0360214, 0.0694630, 0.0464298, -0.0126869, -0.0037262, -0.0008401, 0.0223843, -0.0005775, -0.0002816, -0.0005001, -0.0057539, -0.0471184, -0.0327353, -0.0663711, -0.1279880, 0.0576351, 0.0330379, -0.1129870, -0.2919930, 0.0544826, -0.0133295, 0.1049860, -0.1875480, -0.0183291, -0.0109990, -0.1775060, -0.0000125, -0.0111215, -0.0366339, 0.0773223, 0.0452664, 0.0738452, 0.0360875, 0.0369998, 0.0240618, -0.0012552, 0.0000419, -0.0001605, -0.0073352, -0.0463116, -0.0385386, -0.0976203, -0.0213513, -0.0029332, -0.1588960, 0.0094647, -0.0041713, 0.0334423, -0.0120670, -0.1193350, -0.1532450, -0.1149820, 0.2235740, -0.1562930, 0.0228858, 0.0172371, -0.0398608, -0.0386346, 0.0038011, 0.0027821, -0.0099755, 0.0282647, 0.0043769, -0.0057875, -0.0039030, 0.0001777, -0.0015543, -0.0263043, -0.0124278, -0.1427820, -0.1320820, -0.0957726, -0.1154150, 0.1069110, 0.1022340, 0.0850610, 0.0969757, 0.1200940, -0.2300830, -0.1735410, -0.0777876, -0.1141050, -0.0044669, -0.0473921, -0.0215581, -0.1305230, -0.1255670, -0.0109760, -0.0069073, -0.0039461, -0.0037703, 0.0110227, -0.0000496, -0.0003018, -0.0047254, 0.0202451, -0.0392807, -0.0612130, -0.1040160, -0.0455891, -0.0308313, 0.0388051, 0.0409224, 0.0965757, 0.0343599, 0.0424393, -0.2353710, -0.1698830, -0.0039649, -0.1790790, 0.0374866, -0.0960518, -0.0844338, -0.1015490, -0.1033060, 0.0070564, 0.0417120, 0.0255137, 0.0113482, 0.0043388, -0.0005094, 0.0003674, -0.0112136, -0.0445500, -0.0374877, 0.0109779, 0.1210140, 0.0267400, 0.0917061, -0.0695382, -0.0206438, 0.0209510, 0.0806650, -0.1553250, -0.1363200, -0.1118340, 0.0931358, -0.0953041, -0.0465792, -0.1562750, -0.0465146, -0.0831635, -0.0449896, 0.0574460, 0.0492886, 0.0137831, 0.0106696, -0.0004908, -0.0001211, 0.0002810, -0.0101192, -0.0341137, -0.0699821, 0.1200300, 0.0741975, -0.0153880, -0.0917167, -0.0826925, 0.0531120, -0.2085000, -0.0812777, -0.1269060, 0.0216061, -0.0840878, -0.2517710, -0.1618750, -0.1572030, -0.2018860, 0.0328088, -0.0134273, 0.0364467, 0.1051840, 0.1127500, 0.0216068, 0.0013784, -0.0004315, 0.0005303, -0.0000308, -0.0019692, -0.0101465, -0.0386120, 0.1161360, 0.0959421, -0.0395152, -0.1132990, -0.0868308, -0.1519800, -0.2682740, -0.2020290, -0.0148041, 0.1327560, -0.0538863, -0.1084830, -0.1372050, -0.0215817, 0.0122405, 0.1176180, 0.1210970, 0.1067830, 0.0982309, 0.1089210, 0.0259332, 0.0035715, -0.0000833, 0.0004928, -0.0001665, -0.0012111, -0.0115259, -0.0597901, 0.0817034, 0.0743468, -0.0756773, -0.0429035, -0.0372535, -0.1105120, -0.1175590, 0.1460350, -0.0479305, 0.0022372, 0.0241403, -0.1003970, -0.0778530, 0.0331798, 0.1065670, 0.2022130, 0.0814138, 0.0048119, 0.0472687, 0.0557988, 0.0240474, 0.0117514, 0.0003121, -0.0007313, -0.0000928, -0.0006425, -0.0073665, -0.0638211, -0.0744480, -0.1322120, -0.1095390, -0.1342810, -0.0283894, -0.1031000, 0.1057440, 0.0593422, -0.0247382, 0.1339340, 0.1620490, -0.0858766, 0.0452776, 0.1292790, 0.1853040, 0.1032690, 0.0614147, 0.0208169, 0.0490511, 0.0304337, -0.0005747, -0.0002160, -0.0001375, 0.0003568, -0.0001314, -0.0005728, -0.0013670, -0.0293684, -0.0671483, -0.1431580, -0.1565570, -0.0583440, -0.0536330, -0.2864200, -0.2667200, -0.0603035, -0.0328149, -0.0156739, -0.0340704, -0.0897830, 0.0695359, 0.0445639, -0.0974319, -0.0138242, 0.0409224, 0.0311613, 0.0754883, 0.0302052, -0.0002206, 0.0000508, -0.0000767, -0.0005178, -0.0001214, -0.0002948, 0.0001153, -0.0017846, -0.0169238, -0.0397400, -0.0604930, -0.0452521, -0.0578536, -0.0696375, -0.0582436, -0.1558130, -0.2060260, -0.1627970, -0.1258920, -0.1528550, -0.1159410, -0.1363980, -0.0708708, -0.0408480, -0.0403936, -0.0345008, -0.0050604, -0.0017728, 0.0000873, 0.0003235, -0.0003404, -0.0003975, 0.0001854, 0.0000465, -0.0003051, -0.0000661, -0.0000262, -0.0025358, -0.0125535, -0.0103998, -0.0025883, -0.0075446, -0.0063138, -0.0128138, -0.0158858, -0.0371595, -0.0173698, -0.0166750, -0.0230856, -0.0451698, -0.0092708, -0.0067436, -0.0149084, -0.0214773, -0.0032687, -0.0000656, -0.0003614, 0.0004649, 0.0000898, -0.0002898, 0.0004985, 0.0004500, 0.0000991, -0.0001001, -0.0000764, 0.0003945, 0.0003852, -0.0000609, -0.0002911, 0.0003731, -0.0001509, -0.0005577, -0.0003715, -0.0002080, -0.0001789, -0.0002045, 0.0001405, 0.0002776, 0.0000792, -0.0001888, 0.0003626, -0.0000131, -0.0001765, 0.0001452, 0.0000985, 0.0001559, -0.0002153, 0.0000373, 0.0001194, -0.0000664, 0.0004604, 0.0002712, -0.0002805, -0.0004569, 0.0002540, 0.0005590, -0.0002830, 0.0035120, 0.0130743, 0.0068826, 0.0004265, 0.0030156, 0.0004933, 0.0010410, 0.0011385, 0.0015544, 0.0015235, 0.0006949, -0.0001142, -0.0001499, 0.0004603, 0.0004775, -0.0001445, -0.0000318, 0.0003176, 0.0002731, 0.0003634, 0.0001543, -0.0003181, -0.0004775, -0.0001571, 0.0003951, 0.0010239, -0.0000397, 0.0012571, 0.0233427, 0.0247666, -0.0147067, -0.0006030, 0.0026670, -0.0169077, 0.0160904, 0.0589912, 0.0046108, -0.0412983, 0.0200800, 0.0396126, 0.0134345, 0.0006265, 0.0010781, -0.0000250, 0.0004037, 0.0000018, -0.0001192, 0.0001952, -0.0007746, -0.0015530, -0.0195529, -0.0058880, -0.0102799, -0.0510154, -0.1185240, -0.0458347, -0.0491344, 0.0139900, -0.0853795, -0.0327777, 0.0084458, -0.0327026, -0.0047730, 0.0586492, -0.0630957, 0.0067692, -0.0970776, 0.0424758, 0.1340940, 0.0347830, -0.0299026, -0.0075685, 0.0019966, -0.0007011, -0.0000117, 0.0000376, -0.0028683, -0.0027526, 0.0076358, -0.0082646, -0.0191910, -0.0905323, -0.1079640, -0.0943573, -0.0888104, -0.0234853, -0.0847525, -0.0291617, 0.0155892, -0.2204370, -0.0997102, 0.0426106, -0.1835320, -0.0622527, -0.0533038, -0.1142040, 0.0115237, -0.0417967, -0.2432390, -0.0563279, 0.0143107, -0.0002200, -0.0003785, 0.0000377, 0.0005171, -0.0371056, -0.0110742, -0.0633664, -0.0538562, -0.1472400, 0.0284987, 0.0641704, -0.0451844, -0.1800390, -0.0834155, -0.1260770, 0.0493760, -0.0523161, -0.1465930, 0.0321015, -0.0528913, -0.1632600, -0.1019210, 0.0579374, -0.1011410, -0.0895327, -0.1310870, -0.0237575, 0.0097844, -0.0032303, 0.0000592, -0.0002389, 0.0046994, 0.0313417, 0.0248319, -0.1331540, -0.1271650, -0.0637259, 0.0366695, 0.0463260, -0.0092392, -0.0040572, 0.0281548, 0.0091732, -0.0961097, -0.0382792, -0.0727765, -0.0844064, -0.0771974, 0.0749138, 0.1238340, 0.1301150, -0.0442246, 0.0083824, -0.1623840, -0.1026950, -0.0833154, -0.0112380, -0.0000472, 0.0052225, 0.0109536, 0.0420915, 0.0893222, -0.0778056, -0.0040219, 0.0707304, 0.0125222, 0.0922418, 0.0833327, 0.0111947, -0.1203520, 0.0233588, -0.1172580, 0.0980769, -0.1371760, -0.2962420, 0.0996732, -0.0620581, -0.0750569, 0.0481311, 0.0385116, 0.0124163, -0.1169250, -0.1013820, -0.0248671, -0.0011895, 0.0078952, 0.0086311, 0.0299672, 0.0818970, 0.1480810, -0.0470030, 0.0375862, 0.1772210, 0.0355574, -0.0989067, -0.1723720, -0.1126750, 0.0470393, 0.0881826, 0.0240655, -0.0413238, 0.0657385, 0.0853977, -0.0501391, -0.0308018, -0.1113000, -0.2115950, -0.0543110, -0.0117508, -0.1444950, -0.0699635, 0.0063353, -0.0001402, 0.0003735, 0.0053793, 0.0535331, 0.0862802, 0.1163950, -0.0317268, 0.0147096, -0.0161784, -0.0966031, 0.0513186, -0.0725710, -0.2158090, -0.0539686, 0.0814955, 0.0586487, -0.0324969, -0.0298297, 0.1602940, 0.2491500, 0.2914910, 0.0742768, 0.0022890, -0.1603370, 0.0175500, -0.0624252, -0.0858047, -0.0343889, 0.0005754, 0.0007191, 0.0046892, 0.0399677, 0.0406009, 0.0676647, 0.0025503, -0.0088012, -0.1087880, -0.1520700, -0.0420127, 0.0308703, -0.0961198, -0.0829101, -0.0457532, -0.3039310, -0.1025010, -0.0435463, -0.1130540, 0.1317110, 0.0804804, 0.1578500, 0.1023140, 0.0133341, 0.0931146, -0.0503116, -0.1700160, -0.0568837, -0.0003193, 0.0000370, 0.0100961, 0.0515662, 0.0373175, 0.0227317, 0.1177850, 0.0814387, -0.0156831, -0.0697628, 0.1704880, 0.0078347, -0.0594022, -0.0508035, -0.0149552, -0.1788110, -0.2053210, -0.1330640, -0.2498730, -0.2383570, -0.0177145, -0.0366827, 0.0937395, 0.2395900, 0.2355450, 0.0959072, -0.0134555, -0.0030616, 0.0004939, 0.0003230, 0.0065051, 0.0369470, 0.0567504, 0.0563418, 0.1273050, 0.1679100, 0.0885319, -0.1115640, 0.0381942, -0.2287480, -0.1976800, -0.0806356, -0.1569530, -0.2282000, -0.1287510, -0.0466880, 0.0761571, -0.0412918, -0.0557469, -0.0694355, 0.1224910, 0.2348620, 0.2841040, 0.2299920, 0.0354119, -0.0092980, 0.0006800, 0.0001689, 0.0026392, 0.0339815, 0.0062232, 0.0988822, 0.1819180, 0.3935150, 0.1024190, -0.1499590, -0.0515629, -0.1889800, -0.1288770, -0.2376250, -0.2786580, -0.1344340, -0.0809288, -0.2684640, 0.0003818, 0.0230348, -0.1462030, 0.0400364, 0.0336962, 0.1377710, 0.2634320, 0.1488970, 0.0375816, 0.0033639, 0.0069244, -0.0000244, -0.0034606, 0.0098181, -0.0112483, 0.1437520, 0.4436560, 0.5928920, 0.3636970, 0.3544250, 0.1724560, 0.0515824, -0.0845390, -0.3310110, -0.1129800, -0.1043750, -0.0508192, -0.0681240, 0.1513280, 0.0169892, 0.0487230, -0.0219235, 0.0737655, 0.0687106, -0.0482895, 0.0586460, 0.0501728, 0.0056501, 0.0004356, 0.0007399, -0.0100318, -0.0099404, 0.0028986, 0.0124561, 0.3019450, 0.5429720, 0.8889340, 1.0067400, 0.9083180, 0.5143290, 0.2370330, -0.2697230, -0.2490880, -0.0769323, 0.0605789, 0.0345590, -0.1072520, -0.0873268, -0.0138966, -0.0520459, 0.0494611, -0.0220144, -0.1008810, -0.0378590, 0.0429984, 0.0042083, 0.0038796, 0.0006439, -0.0050777, -0.0199514, -0.0647561, -0.0666409, -0.0169145, 0.1756160, 0.4424700, 0.7480810, 1.1126600, 1.2572400, 1.2486200, 0.7968240, 0.4526670, 0.1057460, 0.0242737, -0.0726976, -0.0300264, -0.0133435, -0.0395217, -0.0703786, -0.0417917, -0.1090100, -0.0517059, -0.1281210, 0.0633089, 0.0166519, 0.0082639, 0.0002817, -0.0016448, -0.0150820, -0.1739500, -0.1011660, -0.0278577, -0.1502390, 0.0137397, 0.0408895, 0.2906480, 0.7777380, 1.0159300, 0.9047670, 0.7603120, 0.3550540, 0.0921223, -0.0833781, -0.1313520, 0.0139719, -0.0891240, -0.0220232, -0.0513911, 0.0513902, -0.0417450, -0.0406124, 0.0953990, 0.0062663, 0.0004816, 0.0008058, -0.0003985, -0.0051747, -0.2955740, -0.1970900, -0.1119340, -0.3576510, -0.2745780, -0.3529820, -0.2249690, -0.2503620, -0.1700730, 0.3089800, 0.4274990, 0.2356210, 0.2170190, 0.1088600, 0.0307979, 0.0598533, -0.0491524, 0.0725023, -0.1382230, 0.0439650, 0.0532417, -0.0901965, 0.0578477, 0.0170213, 0.0000897, -0.0003094, 0.0086955, -0.0150008, -0.2788830, -0.1620020, -0.2141790, -0.2478800, -0.3913730, -0.3115640, -0.1338430, -0.3222640, -0.3770180, -0.1818870, 0.0941920, 0.1599830, 0.2647750, 0.2087260, 0.2404340, 0.0516784, 0.0824794, -0.0503603, -0.1130490, 0.0779940, -0.0879608, -0.1311970, 0.0010759, 0.0052152, 0.0001422, -0.0005821, 0.0001680, 0.0020043, -0.0890619, -0.1184450, -0.2727450, -0.2110380, -0.0320839, -0.2879560, -0.2336620, -0.2096450, -0.2014800, -0.1802100, -0.1053160, 0.0635236, 0.3636210, 0.0288870, 0.1310530, 0.1436810, 0.0993565, 0.0848732, 0.1190320, -0.0624708, -0.1105200, -0.0572975, 0.0157896, 0.0043346, -0.0001365, 0.0009330, -0.0003279, 0.0552219, 0.0727903, -0.0136592, -0.0857696, 0.0208786, -0.1003790, -0.1765950, -0.0437809, -0.1519070, -0.1592220, -0.1457500, -0.2192420, -0.1524780, -0.0432241, 0.1602360, 0.1866100, 0.0907385, 0.1390890, -0.0013288, 0.0464477, -0.0701014, -0.0033641, 0.0272188, 0.0454739, 0.0028100, 0.0001617, -0.0002551, -0.0003352, 0.0503227, 0.0599499, 0.0426480, 0.0532602, 0.1030610, 0.0647904, -0.0000791, 0.0379434, -0.1080110, 0.1135540, 0.1143170, -0.0223199, -0.1798420, 0.0244663, -0.0107512, 0.0515270, 0.0691513, -0.0060224, 0.0786687, 0.0203918, 0.0482132, 0.0370030, 0.0590018, 0.0522737, -0.0004335, 0.0001375, 0.0000173, -0.0002566, -0.0300469, -0.0903577, -0.0573108, -0.1508930, 0.0732497, 0.1245740, 0.1081460, 0.0968285, -0.1339890, -0.1612380, -0.1143940, 0.0468814, 0.0845511, 0.2165780, 0.0520319, 0.0923797, -0.0972616, 0.1238840, 0.1704500, 0.1009840, 0.1220500, 0.0502969, 0.0178969, 0.0311046, -0.0007575, 0.0004398, 0.0000834, -0.0002256, -0.0295092, -0.0651981, -0.0955609, -0.1185680, 0.0047434, -0.1115030, -0.0591175, 0.0407081, 0.0409080, 0.1113710, 0.0738580, 0.0420302, 0.0265534, 0.1118360, -0.0571608, 0.0165061, 0.1770700, 0.2715990, 0.0760082, 0.0805316, 0.0154339, 0.0056265, 0.0166842, 0.0091554, -0.0002193, -0.0005032, -0.0009108, 0.0001405, -0.0049133, 0.0014846, -0.0287308, -0.0608206, 0.0099165, 0.0022635, 0.0060228, -0.0139146, -0.1357490, 0.0374735, 0.0011406, -0.1430370, -0.0413783, -0.0136699, -0.0349933, 0.0271170, 0.1447000, 0.1155280, -0.0211928, -0.0079956, -0.0012061, -0.0078266, -0.0012504, -0.0000279, -0.0001281, -0.0003110, 0.0001206, -0.0000745, -0.0001381, -0.0005101, -0.0107632, -0.0485274, -0.0150230, -0.0011525, 0.0385226, -0.0556109, -0.0984841, -0.0865556, -0.0049773, 0.0708062, -0.0501215, -0.0726626, -0.0555155, -0.0648325, -0.0298188, 0.0377029, 0.0157727, 0.0012251, 0.0073218, 0.0004644, 0.0003041, -0.0000759, 0.0007835, -0.0001249, -0.0000066, 0.0000185, 0.0000610, 0.0002379, -0.0000532, 0.0007304, 0.0014144, 0.0073247, 0.0098842, 0.0120464, 0.0365331, 0.0209590, 0.0254368, 0.0468278, 0.0251925, -0.0410081, 0.0053279, 0.0222692, 0.0167743, 0.0280837, 0.0118577, 0.0007993, 0.0006008, 0.0006005, 0.0002553, -0.0001657, 0.0002048, 0.0001672))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s1,
    done => done_s2,
    start => start_s3,
    ack => ack_s4,
    in_a => in_a_s5,
    out_a => out_a_s6,
    out_offset => out_offset_s7,
    op_argument => op_argument_s8,
    op_result => op_result_s9,
    op_send => op_send_s10,
    op_receive => op_receive_s11
);
interlayer_u70 : interlayer generic map(
    width => 784,
    word_size => 9
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s71,
    done => done_s72,
    start => start_s73,
    ack => ack_s74,
    previous_a => previous_a_s75,
    next_a => next_a_s76
);
bias_op_u12 : bias_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 14, frac => 14)),
    bias_spec => fixed_spec(fixed_spec'(int => 4, frac => 8)),
    biases => reals(reals'( -1.3714500, -0.0223567, -1.1923400, 2.0255800, -0.1508290, -0.3149190, -0.9097960, -0.0888244, -1.4836400, -1.1160700, 2.2643900, -0.5548600, -0.1523720, -0.2297150, -0.1820460, -0.9278840, -1.1400400, -1.1404700, -0.7352880, 0.1199600, -1.5184400, 0.1645080, 1.0912600, -0.9344400, 1.8746300, 1.0565500, 1.4681500, -0.4600640, 1.4199000, -0.6898230, 0.8850680, 1.8038700, -0.5797730, -0.7777570, 1.3278300, 4.4577900, -1.7186700, 1.9009300, -0.3286180, 1.2920700))
) port map(
    input => input_s13,
    offset => offset_s14,
    output => output_s15,
    op_send => op_send_s16,
    op_receive => op_receive_s17
);
sigmoid_op_u18 : sigmoid_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 15, frac => 14)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    step_precision => 2,
    bit_precision => 16
) port map(
    clk => clk,
    input => input_s19,
    output => output_s20,
    op_send => op_send_s21,
    op_receive => op_receive_s22
);
fc_layer_u23 : fc_layer generic map(
    input_width => 40,
    output_width => 40,
    simd_width => 10,
    input_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 3, frac => 5)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 13, frac => 13)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    n_weights => 1600,
    weights_filename => "whatever",
    weight_values => reals(reals'( -0.1980520, -0.5211090, -0.2770550, -0.2810670, 0.4668170, 0.0220185, -0.7085630, 0.1377680, 0.2099480, 0.7104200, 0.7637650, 0.2873910, 0.3529930, 0.5582390, 0.1478920, -0.0020218, 0.0928232, 0.2257610, 0.4544900, -0.2050090, -0.3569980, -0.4647890, 0.0435871, -0.7147170, 0.3696260, -0.0689537, 0.0810571, 0.2590020, -0.1743550, -0.5618960, -0.5237130, 0.4478640, -0.5774280, 0.1477560, 0.4393190, 0.3481740, 0.6176580, 0.0513317, -0.6483990, -0.6544370, -0.1164450, 0.3105830, -1.4780000, 0.7992950, 0.8123100, -0.7679020, 0.4205970, 0.0387268, 0.5250760, 0.3063430, -0.1269130, -0.8490540, -0.0531785, -1.4653900, 0.0282059, -1.2147200, 1.0816200, 0.9578300, -0.0579348, 1.1508800, 0.4503010, 1.0701100, 1.5552400, 0.4260410, -0.2637910, 1.4938600, 1.1400100, -0.5701910, 1.4419600, 0.7355610, 1.3510300, -1.3012400, 0.3000840, 0.1637660, -0.7111510, -0.5860890, 0.4146380, -0.6030600, 0.8870100, -1.2764300, -0.6007220, -0.8382280, 0.1606400, 0.9995420, -0.7705570, -0.5208640, 0.8761600, -0.8085650, 0.2571840, -0.6183150, 0.3009350, 0.8533350, 0.6685460, 0.1097580, 0.1038100, 0.8688460, -0.3532780, -0.9507780, 0.7311190, -0.2622620, 0.9388500, -0.0893599, -0.3753530, 0.2275000, -1.0799800, -0.2919890, -0.5239310, -0.5278620, -0.0912183, -0.5563890, -0.5751370, -1.1565000, 0.8237220, -0.0653934, 0.5042830, -0.0361780, -1.0446800, 0.0667470, 0.0411597, 0.8847980, 2.1622500, -0.7355280, 0.1861030, -0.4346620, -1.1681000, -0.2987250, 1.2279800, -0.4699740, 0.8305360, -0.4901190, -1.1645900, -0.8460070, 0.3495170, -0.6187420, 0.3078050, -0.6387570, -0.5505670, 0.3932630, 0.5726830, 0.5665720, -0.1943710, 0.6999620, -0.0726642, 0.6143770, 1.1395900, 0.4830020, 0.6173370, 1.8153700, 0.5249260, 0.3755050, 0.2466160, -0.4203930, -1.0432200, -1.2672800, -1.4989400, -0.3463770, -0.4007420, 1.2745300, 1.7238300, 0.6963750, 0.9667540, 0.2347750, 0.1401160, -0.1811590, -0.1543850, 0.3935420, -0.1551180, -0.2885570, 0.1261420, -1.1325700, 0.1644180, -1.3838800, -1.0575300, 0.1651000, 0.3106410, 0.4382210, -2.1235800, -0.4632880, -0.1543040, 0.3216070, -0.8043000, -0.2468380, -0.4513580, 1.3515600, 0.0443874, 0.7652210, 0.8666750, 1.0931400, -0.2090030, -0.6175450, 0.4947460, -0.4726080, -0.0685001, -0.8815450, -1.1950200, 0.3954270, -0.2775190, 0.2314580, 0.0749473, 1.7071500, -1.0463200, 0.8856110, 0.2182140, 0.8089880, 0.1263820, 1.0062300, -0.0181958, -0.4585330, 0.1812950, -0.5247180, 0.2131320, -0.7975260, -0.3138820, -0.1441060, -0.9157090, 0.2456680, -0.7969500, -0.2136730, -1.1524000, -0.6283720, 0.1658830, -0.7928180, 0.2717040, 0.2400530, -0.2523470, 0.4305360, 0.8144760, -0.7745100, 0.2011150, -0.2965460, 0.3154280, -0.9331740, 0.8167210, 0.0519024, 0.0718277, 0.3270370, -0.4460630, -0.6629470, -0.9783680, 0.5192720, 0.1947780, -0.7145300, -1.2908800, 0.7028160, 0.0745228, -0.9042660, 1.4273500, 1.2713900, 0.7384840, -1.0439800, -0.0333267, 0.7656920, 0.2778100, -1.1122400, 0.5592620, -0.3301550, -0.0267296, 0.1283920, 1.3985800, 0.7031130, 0.9964460, 0.9471420, -0.0075245, 0.5441310, -1.0082500, -0.0285577, -0.6998960, -0.0731256, 0.8248320, -0.0892768, -0.4487310, -0.8357810, 0.5137860, -0.7972080, -0.2482980, -0.2043660, 1.4047200, -0.8438220, 0.1436170, 0.5259420, -0.2309500, 0.0560263, -0.0881270, 0.2500340, -0.6434320, 0.9507460, 0.4446320, 0.2958020, 0.7868990, 0.0134594, -0.5127350, -0.4218890, 1.2627100, -0.2000300, -1.3457500, -0.1692720, 0.3277570, 0.5896730, -0.3568480, -1.3413600, 0.2146600, -0.3296730, 0.6800240, -0.9321850, 0.9405050, 0.2095020, 0.2510570, -0.3354000, 0.5502560, 0.1790960, -1.3073800, -0.1719650, -0.1085180, 0.0730421, 0.2141150, 0.1273480, 0.5003120, 0.1250450, -0.1533570, 0.0058702, 0.8930100, -1.1980000, 0.1039100, 0.0920572, -1.2895200, -0.3643290, 0.9639540, 0.8537180, 0.6253670, -0.6273240, -0.9319290, 0.9790690, 1.2957100, 0.5565530, -0.2860330, 0.6046010, -0.2238220, -0.6618700, 0.9908330, -0.4057770, 0.1606460, 0.0410816, -0.9500670, -0.0689055, 0.2282190, -0.6068280, -0.9522590, 0.2351310, -0.3948390, 0.2586540, -1.7838300, 0.0573470, -0.2802090, 0.1012430, -0.2883470, 0.3707060, 0.7085740, 0.5779880, 0.8601610, 0.8666920, 1.0509300, -0.8916250, -0.6314650, 0.2655160, -1.1024200, -1.4253900, -0.0030996, -0.3231100, -0.3779060, 0.0076170, -0.3531760, 0.0627841, 0.0629993, 0.9448210, 1.0845500, 1.2865500, -0.6889390, -0.6540440, 1.3892500, 0.9093560, -0.5491830, 0.7479570, -0.6509230, 0.1314970, 0.0915254, 1.0076300, 0.7375480, 1.2398900, 0.0018401, 0.1401620, -0.4582190, 0.3871560, -0.6982350, -0.3144160, -0.8864780, -0.2478170, 0.1211040, 0.6068060, 1.2507300, 0.6558760, -0.2641170, -0.6929530, 0.9075370, 0.2792000, 0.9215050, 0.4268170, -0.3841920, -0.8665750, 1.3008600, -0.1091110, -0.0509400, 0.2971210, 0.6920220, -0.6518630, -0.5759760, -0.4061400, -1.1454200, -1.1030400, -0.6352710, -0.0781023, -0.0955246, -1.3258900, -0.9259210, -0.4061230, 0.0920674, 0.3543930, 0.3522420, 0.2538200, -0.5433240, 0.3203380, 0.6632140, -1.1166500, -0.3223200, 0.7938000, -0.4497340, 1.4783500, -0.8131660, 0.3696420, -0.2845750, 0.4124120, 0.2647480, -0.1918570, -0.3799150, -0.0225519, -0.6465240, -0.3140360, -0.4121920, 1.0678400, -0.2165200, -0.1319590, -0.3594610, 0.0755628, 0.1453890, 1.2550400, -0.1808150, 1.1326000, -0.6897360, -0.6426530, 0.4113340, -0.3335730, -0.9774300, -0.3014410, -0.9336130, -0.3331520, 0.0576964, -0.0984850, -0.1445250, 0.3354090, -0.5893800, 0.0848858, -1.4375300, 0.8275190, -0.4772500, 0.3716670, -0.1828800, 0.6027900, 1.2228400, -0.2209960, 0.0052733, 0.3624880, 0.8338310, -1.0281200, 1.7254500, -1.1724200, 0.5628300, -0.1779570, 0.7012140, -0.9365350, 0.4108080, -0.1950330, -0.0432084, 1.4984400, 0.1613110, -0.8767520, 0.9307460, -0.9473590, 0.4578460, -0.5066030, 0.2784240, 0.9221000, 0.8754230, 0.0176601, -0.9023080, 1.2177000, -0.5379580, -1.9262100, -1.9929200, 0.5986910, -0.8607010, -0.0131784, 1.0871900, -0.4346870, -0.2282130, -0.4201330, 0.3591670, -0.0699300, -1.4504600, 1.0467300, 0.4660680, -0.1963590, 0.0802446, 0.0288120, -0.0416560, -0.3533130, 0.0005140, 0.1645410, 0.0446439, -0.2468880, -0.0827079, -0.0532793, 0.2670730, -0.1783710, -0.5495120, 0.2885010, 0.0369940, -0.0747654, -0.0835998, 0.0263170, -0.1548460, 0.0852267, -0.2068120, -0.2476070, -0.0278734, 0.5102820, -0.4302400, -0.2488750, -0.1257390, 0.2656490, -0.1332600, -0.2900090, 0.0789442, -0.1123980, -0.0014334, -0.2948780, -0.0227319, -0.0871980, -0.0078047, -0.1102510, -0.3812250, -0.0105126, 0.5734420, -1.1312400, 0.6913480, 0.2319320, -0.6995550, -0.4308050, 0.9243000, -0.0664537, 0.8459650, -0.4594130, -1.1537800, 1.0314200, 1.3466000, -0.0781194, -0.3036720, 0.5208940, 0.0800438, -1.0678400, 0.5221310, -0.0932290, 0.6562660, 0.0399286, -0.9319510, 0.1447940, -0.0061389, -0.5807030, -0.9394740, -0.1506640, -0.3824020, 0.7259980, -0.7080990, -0.6188610, -0.0308863, 0.7281370, -0.0057360, 0.4316790, -0.4392120, 0.4895800, 1.0893800, 0.6473610, 0.1307360, 0.6294790, 0.1282900, -0.3861870, 1.3918100, 0.0336208, -0.8395900, 0.3801540, -0.0834514, 0.6300170, -0.3962070, -0.3192310, -0.7617750, -0.4170460, -0.4584310, -0.8166670, 0.1885260, -0.0270564, -1.0637900, 0.8032260, -1.0854800, -0.1935530, -0.1354100, -0.2283220, 0.2379980, 0.4556100, 0.2122040, 0.0429823, -0.0898152, 1.1216600, 1.2232500, 0.2561280, -0.3743840, 1.0148200, -0.6180950, 0.5642810, 0.5922110, -0.5730540, 0.0910908, -0.8822530, 0.4300500, 0.0173331, -1.3354900, 0.6169380, -0.0738066, -0.5380700, -0.4945520, 0.3986190, 0.1126250, 0.4895180, -0.3468200, -1.7100600, -0.0116463, 0.2493800, -0.4164970, 0.2171450, -0.2820720, 0.3998970, -0.0690219, -0.0753090, -1.2652800, -0.0376394, 0.2140020, -1.3029800, 0.9483960, 2.0703100, 2.1117500, 0.7344280, 0.8139960, 0.7675360, -0.0522791, 0.1484080, -0.6454760, 0.7844080, -1.1106500, 0.6005430, 1.0631000, -0.2273750, 0.7106770, -0.5013800, -0.4559460, 1.3679900, -0.7545820, 0.0176462, -1.1608000, 0.2218970, -0.3013480, -0.1685270, -1.2422500, 1.1642900, -0.3313510, -1.3615200, 0.0633742, 1.0807900, -1.0939700, 0.6110380, 1.3437500, 1.4049500, -1.0155900, -1.2770600, -0.5000310, 0.3504740, 1.2745400, -1.1093500, 1.0923800, 0.9631890, 1.0713300, -0.2910440, 0.5250670, 0.1151850, -0.6785670, 0.8630170, 0.0816736, 0.2430380, 0.6594100, -1.0205800, 0.6300060, -0.3156710, -0.1085220, -0.7733560, 0.1672230, -0.3918470, 0.3224730, 0.5473680, -0.1245020, 0.5224870, 0.4623940, -0.5771880, 1.3416300, -1.2110600, 0.0003636, -0.9451130, 0.3050720, -0.2968970, -0.3233050, 0.2687000, -1.8798500, -0.9496990, -0.0329914, -0.3372030, -0.0785311, -0.8428010, -0.2144150, 0.5165620, -0.1019000, 0.4162020, 0.7337540, 0.6645630, -0.0064801, -0.4683130, -0.2748600, -1.3075400, 0.1159140, -0.4978360, -0.7453320, 1.0852800, -0.3568090, 0.1788250, -0.3435870, 1.5521900, -0.0484215, 0.2044140, -0.8494250, -0.3784480, -0.5006990, 0.1522980, 0.2604280, -0.5933740, -0.5709920, 0.7320930, 0.3372540, -0.8629950, -0.3489670, -0.0140045, 0.1742340, -0.7959930, 1.2755500, 1.3077500, 0.2371530, -0.3370690, 0.2268520, 0.4760390, 1.6417300, -0.1984120, 0.1725830, -0.0023754, 0.4122620, 0.4648040, 0.7515420, -0.5912730, -0.1912610, 0.2601340, -0.1883080, -1.1187500, 0.1948640, -1.2345800, 0.0429022, 0.2109870, -0.3045620, -1.1730600, -0.1753680, -0.0560255, 0.0158322, 0.1657200, -0.2276020, -0.0123621, 0.1839860, -0.6183260, -0.0822690, -0.0060930, 0.1217880, -0.1830620, -0.2127160, 0.0834150, -0.1158120, 0.1668740, 0.1516190, -0.1244560, -0.1701380, -0.0453104, 0.2048400, -0.1062630, 0.2416410, 0.1488770, -0.4431560, 0.0411152, 0.1646100, 0.0773262, 0.0288114, -0.1667170, 0.2147510, -0.4253800, 0.3472940, 0.1227750, 0.1629490, -0.0975106, -0.5351410, 0.0255864, -0.0817116, -0.1112400, 0.0005603, -0.0022578, -0.0035227, -0.0053799, -0.0029549, 0.0030085, 0.0021435, -0.0066141, 0.0012212, 0.0010700, 0.0032865, -0.0021162, -0.0056149, 0.0076041, -0.0048746, 0.0000143, 0.0032161, 0.0013504, -0.0034166, -0.0012294, -0.0007563, -0.0063989, -0.0003962, 0.0064854, -0.0089916, -0.0046237, -0.0023477, 0.0036640, -0.0021443, -0.0046865, -0.0021602, -0.0042699, 0.0000080, -0.0009980, 0.0032901, -0.0004464, 0.0006307, -0.0029802, -0.0065969, -0.0035450, -0.0609644, 0.1487510, -0.1738620, -0.0827686, -1.5252800, -0.6889410, -0.2682200, 0.0567552, -1.4633200, 0.5789820, -0.1850760, 0.5759430, -0.0722014, 2.2387500, 0.0439412, 1.9277500, 0.4235970, -0.3847850, 0.4644420, -0.2150100, -0.4134160, 0.3702770, -0.7065320, -0.0494031, -0.1572990, -0.3626240, -0.4146400, -0.1725770, -0.9576200, -0.1634990, -1.1808200, 1.1087600, -0.1039860, 0.3109700, 0.7453910, -0.8706450, 0.0397011, -0.0090144, 0.2686270, 0.2808620, 0.9527860, -0.8947000, -0.6436240, -0.5320770, 0.0875000, -0.9778030, -0.1774680, 0.5592530, -0.0019098, 0.3662310, -0.1292360, 0.1986780, 0.0353152, 0.2019740, 0.7558340, -0.0666211, 0.1347280, 0.0264764, 1.0801800, 0.7399290, -0.5514230, 0.5374680, -0.2763950, -0.1720520, 0.0782692, 0.1078590, -0.1037720, 0.8011160, -0.1378100, 0.2757590, -0.1986540, 0.6802490, -0.8373990, -0.0045777, -0.5282850, 0.0846304, 0.7401370, 0.2077820, 0.7137480, -0.3861090, -0.0891599, 0.1220130, -0.1848430, -0.3193230, -0.1178130, 0.1247620, -0.0057795, 0.1107680, -0.2497660, -0.2176490, 0.4184890, 0.1081170, -0.5929900, 0.5673030, 0.0648421, 0.1494830, -0.2515690, 0.0081364, -0.0030329, 0.0482248, -0.3137540, -0.2303780, -0.2701020, 0.6537170, -0.6125060, -0.4714990, -0.4292550, -0.0027765, -0.3044760, -0.4229400, -0.3695700, 0.1124580, 0.0645554, -0.4411010, 0.0817045, -0.1572010, 0.3583640, -0.3712940, -0.5769160, 0.1746030, 0.0232969, -0.9549160, 0.1948250, -0.6519040, 0.6396660, -1.3093700, -1.5072200, -0.9383370, -0.8015350, 1.4213000, 1.0309500, 1.0198100, -0.2961640, 1.0768200, 1.4455700, 0.7171270, 0.4181540, -0.7712150, 0.9276920, 1.0105300, -0.4532990, -0.2635790, -0.8295580, -0.4632280, -0.3884500, -0.2169300, -0.1553210, 0.6032100, -0.9676360, -0.2253920, 0.5492330, 0.8386800, -0.6956930, 0.7650920, 0.3866490, 0.2571730, -0.8702580, 0.5714340, 0.1063300, -1.1799700, -0.2813970, -0.5374490, -0.1835360, 0.3751710, 0.0854057, 0.0861324, 0.0211031, -0.6389980, 0.8034390, 0.6306610, 0.1962410, -0.7175850, 1.2887800, -1.1320100, 0.0141185, -0.9186520, 0.4299360, 0.4639280, 0.6541840, -0.5694850, 0.6213120, -0.6272370, 1.4546500, -1.5205700, 0.6655460, 0.6596940, 1.2242800, 0.3961130, 0.6295680, -0.1782910, -0.5378360, -0.8494990, -0.4490620, -0.0448028, -0.1408390, 0.1952780, -0.3495580, 0.5222600, -0.1099240, -1.1092700, -0.9724170, 0.1940550, -0.4100240, 0.0327712, 1.1303900, 0.0462761, -0.7984550, 0.8882670, 0.1154670, 0.4911160, 0.2119210, 0.9954740, 0.2515300, 0.2818270, -0.6737420, 0.0569219, 0.4323160, -0.3588790, -0.4044660, -0.1322960, -0.2252700, -0.6010440, -0.7260050, -0.6234920, -0.5284860, 0.0457627, -1.0591700, -1.0780200, -0.6748530, 0.6768170, -0.1383830, 0.2416800, 0.0871363, 1.3642300, 0.4809810, 0.7691750, 0.9835060, -1.0994000, -0.6459240, -0.4139920, 1.2066200, 0.8135430, -1.0685200, -0.3235080, -0.6012340, -0.2093080, 1.2746600, 1.7995600, -0.2662050, -0.9620920, -1.0103200, -0.1516440, -0.6077190, -0.2040150, -0.3445980, -0.0923678, 0.1814450, 0.7006340, 0.1155020, 0.6962460, -0.2077740, 1.4991800, -0.1307520, 1.4731400, -0.2749490, -0.0236635, -0.6396030, -0.3319850, 0.5898220, 0.8051320, -0.4824330, 0.2388650, 0.2569090, -0.8656680, -0.6614210, -0.8653630, 1.7001100, -0.9168040, 1.0449500, 0.8038690, 0.3077560, 0.5158830, -1.1720500, -0.2561510, 0.7423830, -0.7389820, 0.0865786, 1.8295800, -0.0568998, -0.4814030, -0.2236490, 0.7464130, -0.6560690, -0.5698140, 0.0818422, -0.4961410, 0.3282550, 0.3754610, 0.2457640, 1.2495900, -0.2739810, 1.0107700, -0.3867640, 0.7384500, -0.7756450, -0.0618851, -0.8157050, -0.5964960, 0.2890070, 0.8717650, 0.2525000, 0.2767840, 0.2431660, 0.2234460, -0.5172450, -0.2764840, 1.7206000, -1.1331300, 0.5235650, -0.4392500, 0.8674000, -0.2486050, 1.0124400, -1.0062400, 0.2630040, 0.5259990, -0.0072695, -1.1633300, 0.3081110, 0.6302790, -0.5604050, -0.1625690, -0.0367111, -0.6167520, -0.0962039, -0.8252510, 0.9255540, 0.2269340, -0.5121150, -0.0827577, 0.0631274, -0.1325860, 0.2324600, -0.0251018, 0.7407750, -0.4747500, -0.3735590, 0.6035040, -0.1597840, 0.2816110, 0.9025240, 0.3027510, -0.4566140, -0.0289779, 0.2473570, -0.4892950, -1.0665900, 0.8677500, 0.5049120, -0.7617510, -0.4997280, -0.2940920, 1.2608500, -0.7902290, 0.4055380, 0.4037890, 0.0914047, -0.2988990, 0.1393320, -0.0285092, 0.5992800, 1.7849000, 0.3201390, -0.1408830, 0.4080430, -0.4546050, 0.5611650, -0.3779720, 0.1754580, -0.1726730, 1.0110700, -0.3889720, -0.3242470, 0.4269120, -0.5662380, -2.0805600, -1.9560800, -0.5036860, -0.8399710, -0.6480010, -0.2566400, 0.2914330, 0.1550610, -0.3777660, 1.2474900, -0.0303759, -0.6074750, 0.1804220, -1.0084200, -0.2622500, 0.0787127, 0.0915036, 0.6262390, -0.1333490, -0.6351680, 0.3651260, 0.5288390, -0.9077920, -0.1121300, 0.0307775, -0.3628930, -0.2110590, -0.1335340, -0.0120366, -0.3466240, 0.0715740, 0.4617800, -0.1117740, -0.5447360, -0.2434110, 0.4052230, 0.0574273, 0.0701318, 0.4234960, -0.2260680, -0.3424610, -0.2042980, 0.0967820, -0.0605994, 0.1131520, 0.2551460, -0.5832340, 0.2898840, 0.0862301, 0.2407380, -0.3801260, -1.0645900, 0.3732340, 0.2775730, -0.0105988, -0.0329412, 0.4644380, -0.0404095, -0.3206160, -0.0680933, 0.5291330, -0.3005300, 0.5589010, -0.2651150, -0.4661340, 0.5403140, -0.1737560, -0.5601090, 0.6009860, 0.1599520, 0.2992940, -0.8091610, 0.0553563, -0.0598588, -0.2138160, -0.5911010, -0.3245000, -0.2028570, 0.4191490, -0.0486365, -0.2728560, -0.0953254, 0.0286804, -0.3050700, -0.5685170, -0.4976620, 0.6104260, 0.0001974, -0.6143700, -0.0451107, 0.1028630, 0.6244990, -0.2914380, -0.7081870, 0.6194500, 0.1583860, 0.0801587, -0.0425463, -0.5245870, -0.1933610, 0.3066350, -0.2825510, 0.0097523, -0.1600280, 0.4045190, 0.3255660, 0.0739278, -0.0948080, 0.5613370, 0.0963019, -0.0138044, 0.0911233, 0.3394940, 0.1173580, -0.2669740, -0.2966270, -0.2203560, -0.0712249, 0.0804902, 0.3098510, -0.4131000, -0.2947290, 0.1336840, -0.1996280, -0.4127030, -0.4911820, 0.6007780, -0.4026330, -0.5354310, 0.2750510, -0.2971090, 0.2824920, 0.0571376, -0.3849190, -0.0844313, -0.8892930, -0.0854722, -0.3680470, 0.1913330, 0.5109790, -0.0925612, -0.4694650, -0.0426627, -0.3533920, 0.0833602, 1.2700400, 0.1399350, -0.3563830, 0.3163670, 0.3670160, 0.0897592, -0.5719770, 0.2282470, 0.3053130, -0.0545514, -0.1823140, -0.5117180, 0.1403300, -0.1686070, -0.5796830, -0.1872190, 0.0544856, -0.1682160, -0.1193810, -0.8737040, -0.3036980, -0.0046796, 0.2032230, -0.4393250, 0.2642190, 0.1496720, 0.3337400, -0.4006460, -1.1729400, -0.1922600, 0.3567510, 0.9285380, 0.0415246, -0.8289730, 0.8591000, 0.1920080, 0.2286670, 0.9999630, -0.3450640, 0.6283800, -0.7891430, 0.2449800, -0.1908170, -0.9701450, -0.9346680, -1.5130600, 1.9092500, 1.4135200, -0.9041000, 0.3052730, 0.1803830, 0.8862490, 0.5966650, -0.0908334, 0.4211550, -0.7349060, -1.2126300, -0.8291890, 0.2609030, 1.1700000, 0.7518190, 0.4593920, -0.1601250, 0.4379900, 0.2733490, -1.0315100, 1.0412300, -0.6391380, 0.4903720, -1.5813000, -1.1837800, 0.5184990, -0.1319580, 0.7393740, -0.5925480, -0.0649565, 0.0398195, -0.6705560, -0.6745800, 1.1096300, -0.0632442, 0.0692968, 0.2860370, 0.6166680, -0.6166640, 0.8984350, 1.1485800, -0.0223156, -0.7663510, -0.7739390, 0.5172830, -0.2901180, 0.5118620, -1.1372400, -0.1399790, 0.2899200, 0.4198320, -0.7717750, -0.0385518, 0.4222880, -0.0799374, 0.0201187, 0.5488150, 1.4042100, 1.2099100, -0.3154770, -0.7697280, -0.1265600, -0.0695235, -0.7961060, -0.7310590, 0.1557260, 0.0934130, 0.0467298, -0.0893209, 0.4688440, -0.4444030, -0.2433640, -0.3048530, -0.1361470, 1.1718000, 0.0188478, -0.2404040, 0.7508960, 0.0928349, 0.4689350, -0.8315900, 0.0422883, 0.0103650, -0.4540290, -0.2525230, -0.8077970, -0.0217968, 0.0315422, -0.3240590, -0.4065040, 0.0074538, -0.1241580, -0.3436400, -1.0980000, -0.6614650, 0.1816270, 0.1159550, -0.4417400, 0.5002910, 0.2106770, 0.1016510, -0.1542960, -1.2714000, 0.3375510, -0.0626262, -0.1501430, -0.2062520, -0.1129540, 0.0868068, -0.0041567, 0.0762616, -0.4122890, 0.1166200, 0.1725180, 0.2874280, -0.0027961, -0.2966300, 0.2195720, -0.1228050, -0.1004300, 0.1962220, 0.0268307, -0.0971863, 0.0780098, 0.0522100, -0.3068920, 0.0916179, 0.2723740, -0.5238690, -0.0976053, -0.0606113, 0.1608830, 0.0071957, -0.2037490, 0.1227210, -0.3044040, 0.1241020, -0.0122337, 0.2002250, 0.0293732, -0.1065830, -0.1384090, -0.3271420, -0.2366740))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s24,
    done => done_s25,
    start => start_s26,
    ack => ack_s27,
    in_a => in_a_s28,
    out_a => out_a_s29,
    out_offset => out_offset_s30,
    op_argument => op_argument_s31,
    op_result => op_result_s32,
    op_send => op_send_s33,
    op_receive => op_receive_s34
);
interlayer_u94 : interlayer generic map(
    width => 40,
    word_size => 10
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s95,
    done => done_s96,
    start => start_s97,
    ack => ack_s98,
    previous_a => previous_a_s99,
    next_a => next_a_s100
);
bias_op_u35 : bias_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 13, frac => 13)),
    bias_spec => fixed_spec(fixed_spec'(int => 4, frac => 8)),
    biases => reals(reals'( -0.4771390, -2.4595400, -0.3585070, -2.2782600, -1.6620000, -0.5927400, 2.3536400, -1.0658700, 0.6931860, -1.1541800, 0.3591010, 0.6050330, 3.8481900, 1.2168800, 0.5021270, 0.9399850, -4.0082700, -1.5731400, -0.2603360, -0.0182818, -0.4738970, -2.2559500, 2.3056100, -0.2166940, 2.2768000, -0.5589920, -2.3314600, 2.5311700, 1.8106100, 1.5033900, -0.0977505, 3.0942000, 0.6034570, 0.0658099, 0.4124740, 1.7876100, 3.3845500, -0.4803900, 0.5250400, 0.5823320))
) port map(
    input => input_s36,
    offset => offset_s37,
    output => output_s38,
    op_send => op_send_s39,
    op_receive => op_receive_s40
);
sigmoid_op_u41 : sigmoid_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 14, frac => 13)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    step_precision => 2,
    bit_precision => 16
) port map(
    clk => clk,
    input => input_s42,
    output => output_s43,
    op_send => op_send_s44,
    op_receive => op_receive_s45
);
fc_layer_u46 : fc_layer generic map(
    input_width => 40,
    output_width => 10,
    simd_width => 10,
    input_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 4, frac => 4)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 14, frac => 12)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    n_weights => 400,
    weights_filename => "whatever",
    weight_values => reals(reals'( -1.9563100, 1.1958800, 1.9201600, -0.5184080, 1.2445600, 1.5207800, 0.7878220, -0.7625120, -1.6819100, 1.3054900, -1.5287400, -1.9972500, -0.6890370, 0.0823480, -0.5328240, -2.0066100, -1.2962400, 0.6984440, 0.9902370, 0.8611510, 0.8949880, -0.0113621, 1.1751700, -1.6073500, -0.0324651, -1.6048100, -0.4850170, -2.3381400, 0.7417480, -0.9432220, -0.7315970, -0.9052480, 1.1021900, -0.2486710, -0.8049290, -0.1426120, -1.7539600, 1.1555900, 0.0942531, 0.0617613, -1.6021300, -1.5252300, -0.8200200, 2.2186400, 0.2101580, -0.7519420, -1.0950500, 0.7230090, 1.3747000, 0.7629720, 0.7817040, 0.2875430, 1.2705700, -0.6312630, 2.2244600, 0.8949300, -0.0075306, 0.6500750, -0.0146641, -1.5030000, -0.2727840, -0.0242200, 0.8669260, -0.0396165, -1.0667900, -1.4734300, -1.0335500, -0.4992080, 1.2554000, -0.5070150, 1.6346200, -0.6735990, 0.9932760, -1.0806800, -0.5787020, -2.8987300, 1.5919100, 0.4573100, -2.3486000, -0.7269600, 0.2553050, -1.1663000, 2.3371400, -1.9002600, -1.9501700, -0.4708080, 1.7262300, -0.0498612, 1.7588700, 0.9124920, 1.0050600, 0.3632900, 1.1261200, -0.7208020, 1.9421700, -1.7673900, -1.9395200, -2.2463200, 0.6411710, -1.7518000, -0.1617050, -0.0291082, 0.9440480, -0.2055230, -0.4156840, 1.2407000, 0.7142300, 1.0721500, -1.8325900, -0.5341710, -1.5488000, 2.1242400, -0.4030840, -0.5471010, -0.4725330, 0.2892630, -2.2719800, 0.4549900, 0.3140420, -0.3714580, 0.4289130, -2.7635900, -1.5811900, -0.2551020, -1.3107600, -0.5817040, -2.3359900, -0.3325520, -1.8924900, -1.1411500, -1.7089100, -1.0394600, 1.7959200, -0.0312041, -2.0560500, -0.3297190, -2.8887700, 2.1955100, -2.4739900, 1.5247700, -0.2208930, -0.0123532, 1.6791000, -0.6508090, 0.0076537, 1.1798800, -0.3494150, -1.2498600, -1.5849300, -1.9283000, 1.3139400, 2.5833500, 0.3048210, 0.2411400, 0.9512780, 0.3512750, 1.2944700, 0.6522920, 0.7166870, -0.2611480, 0.0969480, 1.6265500, -0.2631810, 2.5827200, 1.1439900, -1.6545100, 0.1454260, -1.7529400, -1.8176300, 1.9960400, 1.0555100, -1.8986900, 2.0441200, -0.2223480, -0.7352320, 0.3033270, 0.9092160, -2.0555000, 0.2818500, 0.3606900, -0.0733809, -0.0190243, -2.1087700, 1.4668600, -0.9541510, 2.0980200, 1.3832400, -1.8907900, -1.8972000, -0.8057860, 1.2141200, -0.8488190, -0.3563520, -1.0385700, -0.6308970, -0.2835770, -0.8948130, -1.7110100, -1.1387100, -0.1816010, -0.2718040, 2.1829900, -0.7749120, -1.8469300, -2.2850200, -1.5434500, 2.0960100, -1.0301600, -0.7527340, 1.6127500, -2.0851000, 0.0856151, -1.7423700, -0.7391900, -0.1895990, 1.3121600, 1.2968400, 0.2417460, -2.9226200, -0.3798320, -0.5744880, -0.0340863, 1.2696400, 1.1872700, -0.5568690, 0.8878520, -0.6027490, 1.4281400, 1.7986300, 2.7599400, -1.5528200, -1.4961600, -1.2153000, -0.6529380, -0.5365030, -0.4280230, 1.9492700, 1.1871900, -1.3192800, -0.5397430, 0.6323090, -1.8743300, -1.1260000, 1.8657600, 1.2703800, -1.1937200, 0.9312790, 1.1360900, 1.6854300, 0.0916286, -1.9187600, 1.7387600, -2.1131200, -0.3732110, -0.6513450, -1.9226900, 1.2375800, 0.8218980, 0.7249830, 0.5880590, -0.8890620, -0.0239126, 0.3154020, 1.0549200, 0.0008329, -1.3662900, 0.2312770, -1.5509100, 1.6512400, -0.4991400, -1.0866900, -1.0970400, -1.2861000, 1.2799300, 0.6573890, 0.1395740, -1.6153400, -1.7994100, 0.5456530, -0.7897760, -0.9532580, -1.0885200, -1.3542800, -1.4325900, 1.1929700, 0.7469510, 1.5074600, -0.9179750, -1.1758700, -1.8765800, 0.6120430, -0.4390660, 1.4193600, 0.1929450, -1.0710200, 1.4062600, -1.9663000, -2.9781900, 0.8010220, -1.6448400, -0.4687260, -0.0136238, -2.3715400, -0.5496280, 0.4971630, -1.9995300, -1.8442000, 0.8236900, 1.6233200, 1.8599600, -0.7914750, 1.2007500, -0.5583130, 0.8776730, -0.3743510, 0.3118870, 1.3630500, -2.2912800, 0.0752995, -0.2932130, 0.0822417, -2.6602600, -1.3209300, -2.1319300, 2.0966300, 1.2491300, -2.6715100, -1.0279100, -1.9802900, 1.5167800, 1.7418500, 1.2904300, -2.3302600, -0.0091999, -1.6801500, 1.6019400, 1.7619500, 0.7816400, 1.3270300, -2.2881200, -0.0585247, -0.0111562, 1.2380900, -0.3967510, 0.0443894, 1.5503600, -1.4554400, 0.8000350, -1.9932300, -1.1821000, -1.2373400, -1.7916600, -0.5997750, 0.8668420, -0.2087760, 0.4892540, -2.7112700, 0.6368730, 0.9853930, -0.3068270, 0.2681510, 1.7418600, -0.1514530, -2.0893800, -1.6302300, 1.6285800, -0.6959410, 2.4168700, -0.2660200, -2.4280900, 1.0930300, -1.1891500, -2.6725400, -0.8160900, -0.2482440, -0.2772240, 1.5503900, 2.2825000, 0.2402140, 0.5204140, -0.0672223, -0.0262678, -2.4703300, -1.5362800, -1.2848000, -2.4551400, 3.2540800, 0.7787210, -2.0351200, -1.5747000, -0.2290730, -1.1395000, -0.2336540, -0.8425040, -0.6582670, -0.1984610, 0.9478290, 1.4506900, -0.2136580, -0.3992250))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s47,
    done => done_s48,
    start => start_s49,
    ack => ack_s50,
    in_a => in_a_s51,
    out_a => out_a_s52,
    out_offset => out_offset_s53,
    op_argument => op_argument_s54,
    op_result => op_result_s55,
    op_send => op_send_s56,
    op_receive => op_receive_s57
);
interlayer_u102 : interlayer generic map(
    width => 40,
    word_size => 10
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s103,
    done => done_s104,
    start => start_s105,
    ack => ack_s106,
    previous_a => previous_a_s107,
    next_a => next_a_s108
);
bias_op_u58 : bias_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 14, frac => 12)),
    bias_spec => fixed_spec(fixed_spec'(int => 4, frac => 8)),
    biases => reals(reals'( -2.6700000, -3.2368500, -4.4698100, -2.1002800, -3.3805300, -5.1092600, -5.0098800, -1.1594900, -4.8861200, -2.0149100))
) port map(
    input => input_s59,
    offset => offset_s60,
    output => output_s61,
    op_send => op_send_s62,
    op_receive => op_receive_s63
);
sigmoid_op_u64 : sigmoid_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 15, frac => 12)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    step_precision => 2,
    bit_precision => 16
) port map(
    clk => clk,
    input => input_s65,
    output => output_s66,
    op_send => op_send_s67,
    op_receive => op_receive_s68
);

previous_a_s99 <= out_a_s6;
ack_s4 <= ack_s98;
done_s96 <= done_s2;
in_a_s5 <= next_a_s76;
start_s3 <= start_s73;
ready_s71 <= ready_s1;
input_s13 <= op_argument_s8;
op_receive_s17 <= op_send_s10;
op_receive_s11 <= op_send_s21;
input_s19 <= output_s15;
op_receive_s22 <= op_send_s16;
offset_s14 <= out_offset_s7;
op_result_s9 <= resize(output_s20, mk(fixed_spec(fixed_spec'(int => 2, frac => 8))));
previous_a_s107 <= out_a_s29;
ack_s27 <= ack_s106;
done_s104 <= done_s25;
in_a_s28 <= next_a_s100;
start_s26 <= start_s97;
ready_s95 <= ready_s24;
input_s36 <= op_argument_s31;
op_receive_s40 <= op_send_s33;
op_receive_s34 <= op_send_s44;
input_s42 <= output_s38;
op_receive_s45 <= op_send_s39;
offset_s37 <= out_offset_s30;
op_result_s32 <= resize(output_s43, mk(fixed_spec(fixed_spec'(int => 2, frac => 8))));
in_a_s51 <= next_a_s108;
start_s49 <= start_s105;
ready_s103 <= ready_s47;
input_s59 <= op_argument_s54;
op_receive_s63 <= op_send_s56;
op_receive_s57 <= op_send_s67;
input_s65 <= output_s61;
op_receive_s68 <= op_send_s62;
offset_s60 <= out_offset_s53;
op_result_s55 <= resize(output_s66, mk(fixed_spec(fixed_spec'(int => 2, frac => 8))));

uPS : ps port map(
    clk => clk,
    rst => rst_sink
);
previous_a_s75 <= to_vec(reals'(0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0156863, 0.2196080, 0.4117650, 0.6078430, 0.7647060, 0.6078430, 0.1921570, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0196078, 0.2274510, 0.6784310, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.8039220, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.1529410, 0.7176470, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9176470, 0.7411760, 0.7411760, 0.1647060, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0156863, 0.5254900, 0.9450980, 0.9960780, 0.9960780, 0.9372550, 0.5254900, 0.1803920, 0.0941176, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.5411760, 0.9960780, 0.9960780, 0.9960780, 0.7176470, 0.1725490, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0156863, 0.5333330, 0.9921570, 0.9960780, 0.9764710, 0.5529410, 0.0352941, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.5333330, 0.9960780, 0.9960780, 0.8745100, 0.3803920, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0156863, 0.5411760, 0.9921570, 0.9960780, 0.9725490, 0.2196080, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.3843140, 0.9960780, 0.9960780, 0.9960780, 0.2392160, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.2313730, 0.9372550, 0.9960780, 0.9764710, 0.3882350, 0.0039216, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0039216, 0.6549020, 0.9960780, 0.9960780, 0.9294120, 0.4156860, 0.0431373, 0.0078431, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0431373, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.5686270, 0.0980392, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.5490200, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.8313730, 0.0901961, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.8235290, 0.9960780, 0.9450980, 0.3333330, 0.3333330, 0.3333330, 0.5882350, 0.9960780, 0.9960780, 0.4588240, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.8235290, 0.9960780, 0.5686270, 0.0000000, 0.0000000, 0.0000000, 0.2000000, 0.9960780, 0.9960780, 0.5843140, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.8235290, 0.9960780, 0.5254900, 0.0000000, 0.0000000, 0.0000000, 0.6745100, 0.9960780, 0.9960780, 0.5843140, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.8235290, 0.9960780, 0.5254900, 0.0000000, 0.0196078, 0.5529410, 0.9921570, 0.9960780, 0.8941180, 0.1215690, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.5450980, 0.9960780, 0.8784310, 0.7450980, 0.7764710, 0.9960780, 0.9960780, 0.9960780, 0.3725490, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0196078, 0.7960780, 0.9960780, 0.9960780, 0.9960780, 0.9960780, 0.9019610, 0.3764710, 0.0039216, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.3960780, 0.7921570, 0.9960780, 0.7960780, 0.6039220, 0.1176470, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000));
done_s72 <= start;
test_out <= shift_range(std_logic_vector(get(out_a_s52, to_integer(sel), mk(fixed_spec(fixed_spec'(int => 2, frac => 8))))), 8)(test_out'range) when to_integer(sel) < 10 else "00000000";
end system;
