library work;
use work.util.all;

package test_data is
    constant inputs : reals := ( 0.5860107, 0.2199555, 0.3368848, 0.3218961, 0.9179956, 0.6033754, 0.5399897, 0.5823666, 0.0162090, 0.8994686, 0.6611612, 0.5382430, 0.5242841, 0.1083759, 0.8681662, 0.2756673, 0.2095378, 0.1805919, 0.6462137, 0.4445746, 0.0349580, 0.2876540, 0.1937561, 0.0250487, 0.6106468, 0.1370069, 0.8056387, 0.2542463, 0.4295769, 0.6056673, 0.5648002, 0.4890641, 0.7336799, 0.9872453, 0.1538092, 0.5360069, 0.0520135, 0.8209977, 0.9606787, 0.1386959, 0.1661568, 0.6394920, 0.5490943, 0.1404275, 0.4945089, 0.1490793, 0.0700357, 0.2994562, 0.2267655, 0.2394792, 0.2421370, 0.8925259, 0.1325165, 0.7671765, 0.7154884, 0.5669313, 0.0614869, 0.6184669, 0.7950070, 0.6419113, 0.1012582, 0.0050820, 0.0629358, 0.9320357, 0.0900054, 0.7161062, 0.4160899, 0.6682278, 0.7648008, 0.6798314, 0.3130169, 0.6855002, 0.0941468, 0.8601665, 0.4227763, 0.7636607, 0.9717141, 0.4133151, 0.6734375, 0.0925695, 0.7827480, 0.8689053, 0.0868421, 0.2113144, 0.4614513, 0.2683381, 0.0189237, 0.8129294, 0.0920045, 0.2497793, 0.9076485, 0.0912745, 0.3754880, 0.7238112, 0.9658751, 0.5697480, 0.5290993, 0.3226925, 0.5731905, 0.9805313, 0.6502176, 0.5278894, 0.3190422, 0.1398481, 0.6731967, 0.7336540, 0.3557988, 0.9413602, 0.1945969, 0.2612163, 0.4968394, 0.0050080, 0.3047606, 0.6755007, 0.4971579, 0.8951367, 0.7640981, 0.8329656, 0.8646787, 0.6864464, 0.4614799, 0.2401798, 0.8246184, 0.9188189, 0.3523014, 0.3653119, 0.0422341, 0.8306378, 0.0129128, 0.8012554, 0.2120021, 0.1908008, 0.6716601, 0.9512079, 0.7306642, 0.1169806, 0.5671442, 0.7634938, 0.2138356, 0.9181540, 0.6741933, 0.2857571, 0.4307768, 0.2453557, 0.2208595, 0.2463724, 0.6246373, 0.6447128, 0.5991296, 0.1206920, 0.0927099, 0.7840294, 0.1120555, 0.7912376, 0.0298562, 0.0152931, 0.1743128, 0.4481288, 0.3588603, 0.3664292, 0.0974833, 0.0703234, 0.9939762, 0.5034342, 0.3974456, 0.5078975, 0.6344699, 0.3638169, 0.5916611, 0.4231628, 0.1017915, 0.4429892, 0.8876334, 0.0462879, 0.9549222, 0.4543056, 0.0170530, 0.7658070, 0.1692385, 0.7317164, 0.0151155, 0.1714130, 0.0050208, 0.5366198, 0.4276013, 0.2847838, 0.1625286, 0.6968008, 0.2812672, 0.6650475, 0.1794232, 0.7982605, 0.6422011, 0.2352478, 0.8235482, 0.3052124, 0.3238148, 0.5826619, 0.0782988, 0.3223106, 0.7195835, 0.0215118, 0.8200900, 0.3510189, 0.4731665, 0.9167078, 0.1064804, 0.6528713, 0.9137408, 0.7976557, 0.8534838, 0.6918045, 0.7691782, 0.0242289, 0.9626058, 0.4340471, 0.5164910, 0.2694424, 0.5712588, 0.7595188, 0.8381850, 0.7848744, 0.1613188, 0.9707255, 0.4160113, 0.3829434, 0.4002666, 0.9324451, 0.6368762, 0.8012865, 0.5943463, 0.2446464, 0.5697906, 0.5364584, 0.4010923, 0.3719889, 0.6844515, 0.3645624, 0.6566033, 0.4963867, 0.6170364, 0.9417784, 0.4096062, 0.4628811, 0.2959286, 0.1397390, 0.3647083, 0.8252571, 0.2321304, 0.9875398, 0.0411054, 0.2443274, 0.3253950, 0.5418811, 0.9872823, 0.3959707, 0.0098824, 0.1812625, 0.9536577, 0.5128194, 0.7776609, 0.8985208, 0.9061467, 0.3012567, 0.2684404, 0.4035019, 0.8762211, 0.6565309, 0.5049178, 0.2054963, 0.4597414, 0.0228230, 0.2387539, 0.1233904, 0.8283603, 0.8962074, 0.7853437, 0.3319063, 0.2110171, 0.6628863, 0.0917831, 0.7550607, 0.0171843, 0.4487637, 0.3047937, 0.3823454, 0.6265713, 0.9541823, 0.5285726, 0.8434232, 0.6456854, 0.1274648, 0.1706516, 0.7963752, 0.1832901, 0.4117934, 0.2133937, 0.1066796, 0.2976359, 0.5936586, 0.7647960, 0.5769983, 0.5301569, 0.2869212, 0.7450713, 0.9420360, 0.3573182, 0.1936529, 0.5552897, 0.1140527, 0.8426961, 0.8085144, 0.0456158, 0.2255645, 0.6063516, 0.4467473, 0.4116545, 0.3234504, 0.1806212, 0.5128584, 0.9954107, 0.0680464, 0.7042908, 0.5918871, 0.1454352, 0.6272480, 0.7491488, 0.8564494, 0.0803186, 0.8239897, 0.0496688, 0.8321391, 0.3556340, 0.5404674, 0.5581803, 0.0280357, 0.1115060, 0.2945191, 0.4742214, 0.2754396, 0.3353042, 0.0666230, 0.0887244, 0.1416313, 0.6828625, 0.2613280, 0.3927453, 0.5665400, 0.7920664, 0.2179889, 0.2553363, 0.2181123, 0.2283985, 0.0988183, 0.8835898, 0.2389295, 0.1801188, 0.4810658, 0.3394827, 0.1096483, 0.2715704, 0.1350871, 0.3993332, 0.8495877, 0.2099426, 0.1116548, 0.2782053, 0.3754126, 0.3166829, 0.6427616, 0.8038535, 0.7698163, 0.1793764, 0.2356065, 0.3517181, 0.1481805, 0.5335596, 0.9813941, 0.0187166, 0.4677723, 0.6514414, 0.7513249, 0.6757983, 0.1829125, 0.1259046, 0.6102354, 0.4732004, 0.5731640, 0.1467460, 0.6905610, 0.2318498, 0.3812276, 0.6162531, 0.4324676, 0.3043549, 0.2527556, 0.7330391, 0.6141240, 0.2074708, 0.8163805, 0.8069598, 0.3631913, 0.4335819, 0.0251073, 0.7822363, 0.6833370, 0.0942472, 0.7240975, 0.3217353, 0.1117711, 0.5726202, 0.1771772, 0.4436223, 0.8560659, 0.9704085, 0.8177052, 0.5521256, 0.6645593, 0.5196027, 0.8796918, 0.0925632, 0.9390178, 0.0243037, 0.9539316, 0.2137452, 0.8104939, 0.0586606, 0.7602617, 0.8197419, 0.6987039, 0.2739910, 0.4459613, 0.9475092, 0.2050576, 0.3475237, 0.6464737, 0.5586295, 0.8012248, 0.9558187, 0.1237816, 0.9830255, 0.2920959, 0.9092430, 0.7406386, 0.1708196, 0.9301795, 0.5063032, 0.4955221, 0.4869707, 0.0670871, 0.5848761, 0.3587823, 0.4005177, 0.2516252, 0.8616748, 0.7863285, 0.5557490, 0.7539249, 0.4296119, 0.4287680, 0.5736971, 0.3947980, 0.2125202, 0.8853927, 0.8028869, 0.6156532, 0.9235449, 0.1298364, 0.7016301, 0.0488320, 0.2302322, 0.6490897, 0.2496751, 0.5256745, 0.8290422, 0.1819630, 0.8347093, 0.3712468, 0.9200826, 0.0008646, 0.0766833, 0.9564567, 0.8768483, 0.0337422, 0.4222452, 0.2745589, 0.5252481, 0.4630091, 0.6485378, 0.6202391, 0.5325065, 0.0863602, 0.5065016, 0.0621051, 0.2192464, 0.3242528, 0.6896726, 0.4357609, 0.3312780, 0.2851983, 0.8378754, 0.5088010, 0.3569825, 0.8065504, 0.9646867, 0.9921419, 0.8941431, 0.2504237, 0.1413694, 0.4269614, 0.7798672, 0.7035556, 0.1154784, 0.4220907, 0.4644042, 0.1878436, 0.9183094, 0.9833135, 0.7265010, 0.0119554, 0.1715161, 0.8983742, 0.0740987, 0.0391549, 0.0845888, 0.7978038, 0.0663861, 0.3726166, 0.5205090, 0.5804579, 0.9662326, 0.4168928, 0.6091329, 0.5147444, 0.3744999, 0.3658940, 0.9240213, 0.8833235, 0.9611757, 0.4108981, 0.1308708, 0.4180323, 0.0308518, 0.3381710, 0.1807837, 0.1688647, 0.8520053, 0.6925982, 0.6225662, 0.7910574, 0.5454284, 0.2672643, 0.5126631, 0.6185154, 0.4854758, 0.8911760, 0.4195637, 0.4967066, 0.7695628, 0.4034992, 0.5548503, 0.3793804, 0.9530918, 0.1146879, 0.7123230, 0.0727818, 0.0520931, 0.7715617, 0.6645843, 0.1369787, 0.4922838, 0.8090654, 0.6167296, 0.2401208, 0.0038112, 0.1001725, 0.6026879, 0.5051876, 0.1690817, 0.4944772, 0.6753215, 0.2769218, 0.6247580, 0.7288515, 0.3710760, 0.7482232, 0.4905551, 0.3843579, 0.8207388, 0.6216635, 0.7853483, 0.0419293, 0.4127998, 0.4088487, 0.4682412, 0.0614430, 0.3153800, 0.2402262, 0.5108655, 0.4548790, 0.4742054, 0.8783450, 0.2589040, 0.2207558, 0.5519774, 0.8409833, 0.2736879, 0.1751206, 0.1170896, 0.0587253, 0.1662411, 0.4083657, 0.1710941, 0.7758415, 0.1158435, 0.2561155, 0.1666438, 0.4572602, 0.3343984, 0.0046089, 0.8775467, 0.4696118, 0.5325157, 0.1153121, 0.3820703, 0.4409217, 0.8928416, 0.5263052, 0.6696783, 0.6512458, 0.9503618, 0.8953151, 0.0791622, 0.2546846, 0.3269650, 0.1721448, 0.1764905, 0.0128337, 0.1370382, 0.0844274, 0.2126241, 0.7215636, 0.1258692, 0.9695107, 0.1013269, 0.1213106, 0.6403988, 0.4321564, 0.8795896, 0.0106714, 0.8240714, 0.1409344, 0.2305189, 0.9196525, 0.2987994, 0.9144566, 0.5363246, 0.9082073, 0.9334676, 0.0966481, 0.1495852, 0.8890441, 0.3611150, 0.5517548, 0.9746879, 0.9540011, 0.3757145, 0.2779290, 0.7806597, 0.6834649, 0.3062818, 0.8312927, 0.6984528, 0.8423700, 0.1694371, 0.3380327, 0.8937273, 0.9407359, 0.2212792, 0.2554684, 0.0403126, 0.1773137, 0.3831992, 0.0553149, 0.8637418, 0.4498773, 0.2967893, 0.0311548, 0.1588024, 0.8382515, 0.5611924, 0.2787798, 0.8797889, 0.7033729, 0.4254720, 0.3657893, 0.7518476, 0.8794571, 0.8860395, 0.4129399, 0.3367164, 0.4857362, 0.7577078, 0.9866832, 0.5322550, 0.5519026, 0.2809709, 0.7416219, 0.5033755, 0.0304798, 0.2745952, 0.3369788, 0.2069580, 0.1044902, 0.9097502, 0.2694050, 0.7358012, 0.5635562, 0.8845974, 0.3293928, 0.8896557, 0.3471427, 0.6474160, 0.2446290, 0.3973835, 0.7313367, 0.2435984, 0.4323796, 0.7616130, 0.0471579, 0.6190651, 0.6221770, 0.3872264, 0.5753417, 0.7384754, 0.9377047, 0.1262462, 0.4308947, 0.7151822, 0.9450018, 0.2496699, 0.6610897, 0.6925008, 0.4226540, 0.8402515, 0.7758078, 0.6812019, 0.4896715, 0.4307816, 0.6406453, 0.0905541, 0.7224796, 0.2148124, 0.7801939, 0.6280407, 0.5883891, 0.0782282, 0.3398616, 0.4115721, 0.2816193, 0.4298613, 0.6864936, 0.3205517, 0.0168760, 0.2093736, 0.5154145, 0.2133401, 0.6211802, 0.3662388, 0.0679313, 0.6341146, 0.2754813, 0.2389911, 0.7191241, 0.4500901, 0.1662083, 0.7436882, 0.2224781, 0.7139475, 0.3422006, 0.1094517, 0.9753904, 0.9828964, 0.4544086 );
    constant weights : reals := ( 2.2779028, 0.4737773, -1.9537905, 1.0490161, -0.1762281, 1.3615162, -0.4837341, 1.9858269, -1.7577574, 1.1540638, -2.8569395, -1.6857722, 1.6538148, 2.5825597, 2.2541005, -2.8486039, -0.7863467, -1.5892754, 0.3346702, 2.0114816, 0.3936245, 1.0985907, -0.3959604, 2.5210604, -0.7023579, -0.5522205, -1.8895310, -1.3583465, -0.8815659, -2.9506116, 0.8154919, -1.3926852, -2.6760174, 2.7169499, -0.2702609, 2.6584253, 2.4835975, -1.2485674, 2.8372248, 0.6682770, -2.0492260, 1.3641864, 2.3147348, -0.9828280, -1.4552595, -2.5866038, 1.3243875, -2.8663436, 1.4502279, 0.6107989, -2.6927444, -2.7541332, 1.6729054, 0.9854830, 0.3053400, -0.8121092, 1.0152177, 2.5674126, -1.1710885, 0.9180814, -2.2923390, -1.5771671, 0.7644643, -0.1305639, -2.9476435, 1.1853518, -0.2745247, -0.7573082, 0.0406655, 0.4745180, 1.2797387, -0.9146734, -2.6167326, 0.9841840, 1.2008909, -2.5745519, 1.8465690, -1.2477594, -0.8257353, -2.1529116, 0.6333326, 1.5776152, 1.7806423, 2.9494489, -1.3783474, 0.1309367, -2.7538698, 1.1867860, -0.4580025, 1.9417276, -2.7472623, -1.4578771, -0.9220389, 1.7695745, 1.7953972, -0.3619993, 2.7882425, 1.1522876, 1.9561973, -2.6845571, -1.3021694, 2.7697345, 2.7316648, -0.5500277, -0.1084452, 0.3279131, -0.7797791, -2.8098113, -2.6646275, -0.1774489, -2.0913689, 0.0532960, 0.6362620, 2.0075477, -0.4702305, -0.0300334, 1.7691988, 1.9670738, 2.5171759, 2.5207138, -0.6436784, 1.2806244, 0.6802414, 1.4667353, 0.2882208, 0.8502488, 2.2182401, -2.0451211, 2.3341758, 2.1646687, -0.5736463, 2.1859913, 2.7486109, -2.3643804, 2.9098164, -0.7571274, 0.3706965, 0.7172666, -1.0050114, -2.9047726, -2.3122450, 1.3168063, -1.1223610, -1.0323854, 0.4882202, -1.6571812, 1.7966587, -2.0929329, -0.2214641, 0.0297973, 0.3421307, 2.2246268, 0.3163441, 1.5692532, 2.2263677, 0.6167405, -2.7341243, -1.0042222, -2.0959231, -2.5079107, -1.7374597, -0.4314007, 2.5925069, 0.9273748, -2.9652671, -1.8763547, 1.0277310, 1.9630484, -0.6414145, -2.7222067, -1.2166261, -1.7583865, -0.6347550, 0.8706183, -1.1885001, -2.3734086, -2.4410239, -1.2364207, -2.1391623, 0.6417424, 1.1960390, 2.4299180, 1.0509422, 2.5494552, 2.6794006, -0.5051708, -2.2709465, 1.6224251, -0.9338322, 0.5458922, -1.5719258, 0.1940116, 2.3654501, 2.9536920, -0.4905545, -0.2010266, 0.7802982, -1.3414798, -0.4686955, 2.2365787, 2.1756207, 1.5301857, 1.4922902, -2.1389784, -0.0655697, 1.9402862, -2.4538465, -0.4083320, 1.0185465, -0.3323612, 0.5687693, 2.4756081, -0.1794539, 2.3806367, 0.4616833, 1.8458268, -2.2150003, -2.6373314, 2.8696187, -0.3993478, 1.8148522, 2.0162729, 1.0215236, 0.8000315, -0.3975319, 0.1249378, -0.2606096, 0.9988528, 2.2056127, 2.8404060, -2.2799863, 0.3812867, 1.5410095, -0.4893893, 1.8402779, 1.1331092, -2.5175565, 0.6024369, 0.4923395, -0.3056072, 0.6079681, 2.1660915, 0.2181380, -1.2923334, -2.1300455, 0.5409435, -2.8678456, -2.7014763, -2.7804456, 2.2323259, -0.0691828, -0.9107975, 1.6467089, -2.3793411, -2.6612614, -0.8026324, 1.5858621, 2.6904207, 0.9693994, 0.4375685, -1.9334688, -1.6340018, -0.4910066, -2.4761057, -1.0506173, 2.8631394, -0.8395516, -0.9836054, 0.1194301, -2.7581851, -0.3649766, 2.5589754, 0.6797431, 2.1487158, -0.9429275, 1.0819448, -2.2933469, 2.9709521, 0.1900417, -1.4457577, 0.2853173, -1.6565571, -2.6027787, 0.5203940, -1.8793190, -2.3222240, -1.6631776, 0.0806745, 1.4577680, 2.7592179, 1.3330337, 0.8325779, 0.2815843, -2.9224191, -2.2891097, -2.4852209, -0.6798841, 2.6426588, 0.0087216, 0.7874192, -2.3574467, 0.0297743, 2.7769862, 0.1372073, 2.9720962, 0.3076015, -2.0355675, -0.6173804, 1.2071123, -1.0082900, -1.1916894, 2.0475599, -2.7971882, 2.1802879, 2.2098687, 1.8628088, -0.1639807, 0.0675291, -0.3363447, 0.5237377, 1.6262961, 1.6753777, -1.0836668, 1.6857290, 0.9897128, -1.7884189, 0.8078983, 1.2908615, 0.9539245, 1.0106096, -1.2503296, 2.7494697, 2.9847084, 2.1595652, -2.2506976, 2.5481338, 2.9294549, -2.3615513, -2.0372241, -2.5909605, 2.6873631, 0.8603269, 1.2720605, 2.8535511, 0.5406488, 0.1851766, -0.3831216, -0.4978130, -0.5718257, 2.9014845, -2.1195579, -1.9733620, 0.8231128, -2.3973263, 0.3518615, 2.8356543, 1.8086437, 2.7654481, 2.1602044, -2.1306159, -1.0354527, 0.4183871, 0.1122756, -0.3303173, 0.1823544, -1.6664460, 0.0782990, 1.4370612, -1.8412720, -1.5444843, 2.2081930, -2.0806972, -2.4501794, -0.0000105, -1.5290412, 2.7730612, 1.8890158, -2.6912006, 1.0164269, -0.4704674, -1.2490560, -1.6625719, -0.8480458, -2.5816200, -1.8940700, 2.4816175, 1.8302174, 0.8508357, -1.1179295, -1.6846443, 1.7738058, 1.9968041, -1.3534215, 1.9158502, 0.3981609, -1.3247888, 1.9881345, 1.8811504, 2.5063516, 1.3412614, -1.4222976, 2.1355279, 1.1699984, 2.6241585, 1.3411218, -1.8019014, 1.2734760, -2.2786646, -2.8396177, -2.3432579, -0.0721861, -0.3609209, -1.9481057, -0.5165749, -2.5557954, -2.6419486, -1.8738522, -2.3356324, -0.3816157, 2.8033481, -2.7182556, 2.0497549, -2.0379079, 0.4027124, 2.7781337, -1.5423648, -0.1729184, -1.1289950, -1.5420580, 1.5571984, -1.7494018, -0.5949698, 0.1873913, -2.6744836, 1.7163522, 1.7040504, -2.5306129, -2.9885920, 0.7734708, -1.5347781, -2.9114755, 2.2699453, -2.5716728, -2.4884480, -1.1691795, 2.3024459, 0.7388135, 2.8088312, -0.7165262, 2.3054988, 1.4364895, 1.2228661, -1.5544069, -2.1464208, -0.5367780, -0.1634480, -2.2807969, 1.9343593, 2.1997535, 0.2048217, 0.1816403, 1.1687209, 1.2741765, -1.9194967, -0.1076471, -2.6384881, 0.2667214, 1.0900848, -1.2577911, 2.1053824, -0.0112827, -2.4873764, -2.4790887, 2.8825657, 2.1516656, -2.1780694, -1.6527722, 1.8425596, -2.8283579, -1.9861135, -2.2996725, 0.1882647, -0.7565880, -2.2660377, -0.1856972, -2.4338185, 0.5318162, 2.6544601, -0.0841052, -0.4915025, 2.5133506, 2.1863693, -2.5680069, 2.2514898, 0.5118837, -2.3013544, 1.1973956, 1.5258766, 0.4849521, 1.8069937, 2.5511226, 2.8014794, 0.7617039, -2.2892594, 2.7786087, -1.9708892, 2.6389096, -2.9066258, -1.6916066, -1.2443394, -0.8869042, 0.8581460, 0.5475532, -0.8765017, -1.3001087, -1.1772975, -1.6444654, -2.1469080, -1.4406403, -2.7242796, 2.9476512, -1.8471528, 1.9714420, 1.7823916, -0.5560094, -1.1357463, 1.4246147, -2.4605969, 0.6875278, -0.1992626, -2.3196047, 0.1671797, 0.3829740, 0.8907254, -1.3580381, -0.1295449, -2.8699035, -1.0428688, -0.0595525, 1.9038768, -0.7020802, 1.1220794, -0.8813711, -0.9376785, -2.4299965, 2.8345641, -0.3419173, -0.3015299, 1.4368305, 2.2855463, 1.6562434, 1.3570212, 1.1506522, 0.7348157, 2.6535951, -0.2003452, 2.9435844, -1.9288753, -1.2494335, 0.6242472, 1.3165129, 1.7855581, -1.3456458, -0.7521440, 0.1336541, 2.1016119, -2.8079511, -0.8508737, 1.7764365, -0.7193142, -1.3217929, 0.8123389, 1.6091770, 0.2222221, -1.5531611, -0.9147335, -0.9263163, 2.0140278, -2.1940285, 1.5464853, 2.6597376, 2.3000047, -2.7827564, -1.6400824, 1.9969001, -1.4437983, 0.7973245, 1.4554733, 2.7981366, -1.8782921, 0.1813791, -1.5692203, -0.2296621, -2.9377007, 2.2679417, -0.2961495, 2.3502806, 1.7727515, -2.3495984, 0.5486565, -1.5496063, 2.1253244, 1.7873356, -1.6961554, -2.2968213, -1.9883245, 2.8081369, -2.9814495, 2.2740916, -0.1635340, 2.2302124, -2.6486836, -0.9573110, 2.1518274, 0.9846637, 2.7936657, -2.7978216, -0.7027860, -1.9569989, -2.3589629, -2.8704608, -0.7951451, 0.3337136, 0.1791296, -2.3270748, 0.8173646, 2.4343857, 1.6260003, -1.2328466, -2.4244101, -0.5609110, 1.9685013, 0.5916892, 1.6581050, 0.5428573, -1.9293771, -0.8003066, 1.2983126, -0.9822787, 1.7084876, 1.5640488, 2.4360353, 1.3838402, 1.9107948, -1.3959417, -0.5114618, -1.4635549, 2.0421386, -1.2745115, 1.4699880, -0.7263092, 2.3561575, -1.1351092, 0.5261703, 0.5906741, -1.0153541, -0.8979315, -0.5017728, -2.6779109, -2.5887168, -2.3515461, 2.7446092, 1.1038287, -1.0055453, -1.7075784, -1.8550728, -1.5668090, -2.4956066, -1.1885192, 1.5019836, -0.8044511, 2.0872021, -1.4970918, 2.1719596, 2.0620982, -2.0668996, 1.6237990, 0.2523908, -0.4463525, -0.9810314, 0.9705517, -1.5768778, 2.9584986, -1.7382313, 1.1480713, -2.3927549, -0.2761464, -2.0204560, 2.3557952, -0.0540983, -2.1466167, -0.8663708, -0.1567485, 1.5066167, -2.1244243, -1.0857215, 0.8573998, -0.4288160, -2.5666831, 1.0144786, 0.6210781, -2.8343147, 1.0361040, -0.6877903, 2.4717696, -0.2757326, -0.1674980, 1.4007533, -1.0518757, 0.9297839, 2.1388114, 0.8021020, -1.0346575, 1.7006787, -2.1063387, -2.5025537, 2.6835798, 0.8232425, 1.5915007, 2.2996885, -2.7492247, 2.6801654, 2.9917587, 1.9303135, -0.7401684, -1.7335236, 2.5204846, 2.2837656, -1.5179057, -0.4037160, 0.7501016, -2.5159950, 2.9671973, 1.6087249, -2.0956914, -2.7532768, -1.7679019, 2.3480734, 1.3904166, 0.6652145, 2.8494977, -2.0540961, 1.7329807, 2.6775943, -0.0201217, 0.0853684, -1.8599968, -1.5987834, 0.2007210, -2.8372557, 2.7693375, -0.8243489, 1.1951557, 2.2105235, -2.3857197, 2.7034529, -2.3901934, -0.8381375, 1.6318612, -0.3052051, 1.3267470, 0.5910698, 1.6735574, -0.9082194, 2.0383474, -2.7401578, -2.0533466, -0.2682449, -1.4525852, 0.3634116, 1.0807889, 1.9853310, 0.7591772, 1.3878745, -2.1174974, -0.7817984, 2.8884926, 1.0541324, -2.4406464, -2.6022695, 1.2550883, -2.3123381, -1.6429592, -1.6259357, -0.1250918, -0.5296480, 0.7941677, 2.7153502, 0.1611803, 2.5155896, 0.8609876, 2.6846090, 2.0261506, 2.1139774, 0.0577920, 0.2742531, 2.7997099, -1.3899875, -0.0998130, 0.8887210, -1.1637842, 1.8411572, 2.5505568, 2.6705701, -1.0902631, 1.8090345, -1.1994832, 1.6267029, -2.9711801, -1.6248361, 1.0318974, 2.8605161, -0.9660477, -0.5289601, 2.5681225, 2.3696684, -2.5933211, -1.3229690, -0.8978456, 0.1331384, -1.3765736, 1.3593822, -0.7956326, -1.6953630, -1.9506242, -0.4701041, -1.4750923, 1.4141004, 1.9891120, 1.5348499, -1.3780878, -0.3188978, -2.5158847, 0.0495568, 2.7145500, -1.2090502, -2.8974263, 1.9770473, -0.7885613, -2.4902925, -0.9131395, 0.0774583, -0.0918573, 0.4761627, -2.4829339, -2.9464738, -1.5994459, 1.0465110, -1.5059680, -2.7830070, -1.4715798, 2.6313877, 0.8118585, -1.1303511, 0.3986825, -2.6557880, -1.4143521, -0.8125876, 0.3156000, 0.5170833, 0.2349594, -2.2567804, -2.0195414, -2.7665028, -1.8447528, 1.0819638, -0.6827261, -0.2138550, 0.2582700, 0.7752851, 0.5483828, 2.8887351, -1.1304615, -0.5864838, -2.4605215, 2.5011619, 2.2177252, 2.9470462, -1.1431999, -1.1160747, 2.2316511, 1.8146330, 2.7082517, 1.4122531, 0.5781921, -0.3731240, 0.3572843, -0.4277312, -0.5823562, 0.6473866, 2.9424752, -0.2331035, 1.0699101, -0.8209967, 0.9581720, -0.2941102, -2.5560696, 0.8843951, 1.7388558, 2.8692927, 2.0453959, -0.5208413, -1.6524618, -0.0007978, -2.7956264, 0.2076629, -1.5504190, -2.9875376, 2.3384293, 2.3902147, 1.7902946, -2.9293789, -0.6587053, -2.9173302, 2.4808726, 1.1240140, -2.1227113, -1.2406217, 2.0237895, -0.6052272, 0.2200225, 1.5278962, 0.5777225, 0.4618612, -0.9899148, -1.6797204, -2.8116201, 0.3609031, -1.6574601, -1.2644644, 2.2926578, 0.7217248, 1.7119984, -1.5540372, 1.7168227, 1.8552512, 2.1936989, 2.9747448, -0.8716441, -2.6460131, -0.1808933, 2.5909037, -0.7521202, -2.6021355, -1.2787137, -1.8301056, -0.1227138, 1.2948586, -2.6671080, -0.0419284, 1.1372065, 2.8449399, -2.7062852, 1.0470322, -0.7999794, 0.0993468, -0.5064156, 0.2421364, -1.0520178, -0.2911816, 2.8784586, 1.4383622, 2.2417228, -2.4656488, 2.5224768, -1.9682780, 1.0891290, -2.2257868, -2.5572522, -2.3575294, -1.8955177, -0.8178454, 2.6055276, -2.1956357, 0.3297573, 2.2955775, -2.1479255, 1.0389034, 1.9560615, 2.7358116, 0.1509263, 1.2137070, 2.1585946, 2.0691482, 1.6793293, -0.9125759, 2.7436480, -0.3337252, 1.8949090, -0.1643261, 0.8987791, -1.8986892, 0.9672810, 1.0260392, -1.1559599, 0.6620582, -2.6631623, -0.7385927, -2.5832066, -1.8961895, 0.7887230, -1.7521725, 0.4251573, 1.3286762, 2.3283667, 1.1745794, 2.6278952, -2.3459503, 1.8223885, -1.2794735, -0.8566010, -1.2295819, 0.3013576, -1.0444421, -2.1628957, -2.5626302, 0.7982909, -1.6836906, -1.5472122, -2.5612155, 2.3446432, 2.8816382, 1.9825320, -0.9651391, 0.7236545, -1.9360494, 0.1053318, 2.0505529, 0.9600224, -0.4235746, 0.0406115, 2.7153780, -1.3400749, -2.2364412, -1.4073828, -1.6201852, -1.0424380, 0.4704615, -1.6664899, 0.8900661, 1.0757534, -0.8052629, 1.5824455, -0.5094669, -0.4131436, 2.0088913, 0.2835037, 2.4668120, -1.7212601, -1.5972186, -1.8158976, -0.8994815, 2.7861991, 0.6556144, 0.5379630, -2.8535631, -1.4246616, 1.5496135, -2.4260204, -0.3250671, 0.4245893, 0.2397881, 0.7922366, -2.2778288, -1.2159167, 0.8061846, -2.1420146, 2.8925355, 1.1658303, 2.3330553, -1.0308709, -0.3322153, 1.5057756, -1.9026943, -1.3347300, 0.2609736, -0.9352206, 1.1155215, 2.8862880, -2.1404182, 1.9773782, -0.4433616, 2.5732290, 0.2916657, -0.3048158, -0.3608064, -1.7991142, 0.1561339, -0.3361723, 0.1679340, 2.1241143, 1.3820732, -1.4949801, 2.5919802, 2.5561583, -2.4335902, 0.5014339, 2.6572705, -1.4698391, -1.7978377, -1.8974546, 0.2628055, 0.8753386, -0.7647799, 0.0441799, -1.4668669, 2.1168959, -0.1459715, 0.3947025, 0.3649271, -0.1499150, 1.9495598, 1.1932113, 2.9191719, 2.5998698, 0.9570932, -0.1722945, 2.5467213, 1.2276151, 2.5687302, -2.1502357, 0.7333064, 1.5262913, 0.6382402, -1.3647825, 1.9828064, 0.8225844, 2.4101582, 1.6535673, -2.3027097, -2.4596793, 2.5759878, -2.1754959, -0.9607558, 0.4921109, 2.4148934, -1.0933553, 2.4971042, 0.0570257, 2.5786142, -2.0266584, 0.6638212, -1.1960538, -0.2961871, 1.8168365, 0.7906398, 0.8626955, 0.0030475, -2.8632920, -2.2252291, 1.4574414, 1.1459414, 1.8223285, -2.2733290, -1.9383135, 1.4043457, 2.6778304, 2.3170400, -0.9231192, -0.2849615, -0.4488993, -0.1961207, -0.5299571, 2.6540467, 2.9868294, -0.4918178, -0.3630171, -2.0150678, -0.0863734, -1.0632449, 1.1003289, -1.7410770, 2.6191523, -2.0555378, -0.1184993, 1.2937484, -1.0603323, 0.2318636, -0.0738532, 2.7776565, 2.6808250, 0.9458553, 2.0931179, 1.6444299, -0.3213381, -1.6046804, 1.3541409, -1.0805295, -2.4630258, -1.1972528, 1.3040460, 2.8808587, 2.3768931, 2.2439328, -0.7847123, -1.3350205, -2.6794799, 2.6508672, 2.3944232, -0.4854233, -1.2684931, 2.2878390, 2.2124164, -1.3580131, -1.2058194, 0.5868537, 0.4337891, 2.7439769, 2.4005670, 0.6247731, 1.5858495, 2.8627051, -0.8427442, 2.5628566, 0.6683446, 0.4603859, -1.2374174, 0.6113833, -0.4088221, 2.1203398, 0.6245556, 1.7758619, 0.4750708, 1.3891622, 1.9628417, -1.2104216, 1.7853383, 1.1065555, -2.6341228, 2.6269552, -0.6434416, -1.1756654, -1.6237041, 0.3253034, 2.3231512, -1.7765742, 2.4932039, -2.7978099, -2.8502027, 0.0476503, 2.6275537, 2.0391364, -2.2621725, 1.1492860, 2.7442749, 1.0336901, -1.3192710, 2.6072727, 2.1128829, 2.1996857, -0.0261328, 0.0579712, -1.8378064, 1.7336201, -1.6747061, 2.5182938, -2.2587322, 0.4795094, 1.8708297, 2.3337490, -2.5602887, -1.5406214, 2.0450105, 1.4265992, -1.8849502, -2.1812443, 2.5696580, 1.1627375, -1.5449315, -0.7282899, 2.4244803, 2.8259415, 1.8758626, 1.6229908, -0.5994261, 1.9543903, 2.3791507, -1.8898582, -0.6991005, -0.2458763, -2.1047116, -2.0526577, 1.3214559, 1.8119146, -0.4893705, 0.5090688, -2.0968979, 0.7405759, -1.2791992, 2.2125185, -2.3509721, -0.2976646, -2.4836710, 1.8825865, 2.8168320, 1.8668127, -2.7217556, 1.2046704, -2.6239512, -2.8391492, 1.7633795, -2.2809413, -0.3574871, 2.5237519, 0.8988340, 1.9661971, 1.4476533, -0.6789082, 1.4464420, 2.9758015, 1.4153629, -1.9408349, -1.7305013, -0.3367840, -0.4051037, 2.6474145, 2.4026469, -1.7167544, -1.6954846, -1.2933112, 0.2498030, 1.6652976, 2.3819265, 0.7224736, -0.8029460, -2.6050010, -2.1479779, -1.7334242, 2.3343467, 1.5683475, -0.3489372, -1.0944333, 1.2593666, -2.1613569, 0.9295559, 0.6395646, 2.4357253, 1.8952782, -0.9458258, 0.2762992, 0.4993481, 1.1265848, -0.7329691, 2.1310845, 0.6461385, 0.9884610, 1.6702618, 0.7191974, 2.8527542, -1.3667609, 2.2185441, 2.0526142, -2.7611429, 0.5427735, 0.3081114, -2.5820594, -2.5292394, 2.6450506, -1.3636344, -2.2309220, 1.8831083, -0.9865224, 2.3861974, -1.2720612, 0.4076305, 1.7517420, -1.6790820, 1.2022086, -1.8658141, 1.4684103, 1.0105937, -0.3855040, -2.0261340, -1.6167352, 1.6441903, -1.8711388, -0.9683311, -0.9272961, 1.6053545, -2.8887638, 0.6780440, -1.7609338, 2.3410924, -2.7505533, -0.9971780, -1.0273176, 2.4825861, -2.6730398, 0.3509188, 2.6840220, -2.3497990, -0.1439248, 0.1372813, 0.9385852, -1.5371401, 2.7005892, 1.8090787, -2.9217694, -2.6679431, 1.2989395, -0.6492534, 1.7397053, -2.4335319, 1.3957234, -0.1997998, -1.8667177, -0.6188009, -0.7809848, -1.6866300, -2.6156083, 2.7007074, -0.3363399, 2.5662312, -1.0828648, 1.5700397, 1.4471669, -2.2387788, -0.2479913, 1.5667690, -0.2408105, 0.9568473, 1.9730303, -1.6547432, -0.5871321, 2.9179944, 2.9891329, 1.1954475, 2.0777900, 0.9738475, -0.0107527, 1.8618814, -1.6304357, -1.5351620, -0.5236547, -0.3738616, 0.1290480, 0.3075027, 2.9075856, 1.4911493, -1.4039902, -0.9631187, -0.0203960, -1.2278973, -1.2845758, -0.1464515, -2.5700785, 1.3283445, -2.9202007, -0.1303023, -2.4605516, -1.1469183, -1.7121229, 1.8215694, -0.3920353, 1.0613400, -2.4418991, 0.5353782, -0.2786034, -0.6402602, -0.4780089, -2.9336067, 2.2585357, -2.0808332, -0.3974529, 1.4477296, 1.5191022, -2.9195771, 2.8713940, -0.1582947, 0.0025742, 0.0484708, 2.2600389, -1.0895207, 1.3490251, 0.8631122, -2.4575268, -0.4958819, 2.1096286, 1.1112305, -2.8896835, 0.6207063, -0.1639300, -0.7508929, -1.8431981, -2.1389639, 0.9906908, -1.4484175, -1.6509661, -2.9138954, -0.0754470, 2.3838977, 1.3725635, -1.0674397, -1.6693003, 0.3271014, 2.9553508, -2.3524724, -2.9655278, -2.0359500, 2.8909127, -0.6147647, 2.8845996, -1.6507578, -0.4142571, -1.0659385, 2.7477371, -1.8494626, 1.0969453, -1.2634041, 0.2495154, 2.0193714, -1.2327719, -0.2021871, -0.9216927, -2.2811227, -0.0306740, -1.6365718, 1.7109662, 0.5868483, -2.1285444, 1.7241643, 1.3781566, -1.0834839, -2.5600936, 0.4028524, -0.5869837, -1.2576199, 2.2508244, -1.3637384, 1.2230255, -2.5138808, -2.2309880, 2.8217128, -1.2264641, 0.1823460, 0.1552094, 1.0272453, 2.2493505, 1.2880581, 1.0845555, 2.5367965, -1.6769802, -1.7486601, -0.9323736, -1.5216426, -1.9962525, 1.5387276, 0.3286751, 0.6016626, 1.9670387, 2.7811727, -2.1019674, 2.7558665, -2.5191711, 0.8972439, -0.0140469, 0.3340023, 1.0940893, 0.7487358, 2.5440893, 1.9441765, -2.5747545, 0.9794785, 0.4685901, -1.1002450, 1.2958207, 1.6515451, -0.9206224, 1.5803405, -1.1380253, 0.9263029, -0.7918731, 0.9566031, -1.5779569, 1.1754947, 2.1532478, 0.3798186, -2.2908239, 1.5789238, -1.2239851, -2.4209045, -2.1020184, 1.7924201, -0.8587985, 1.9144771, 2.3834579, -1.8799594, -1.7098651, -0.5296090, -1.8174715, 2.6080011, 0.4957207, 1.0659190, -0.6885419, -0.2423582, 0.0894142, -0.6912925, -2.1587318, -2.9647535, 2.3326859, 0.2982092, -1.2225655, 2.0331424, -1.6414874, 2.1706369, -1.2501645, -2.4817599, 0.7784868, 0.3171897, -2.4133862, -2.7753313, 2.8578987, -1.5928401, 2.8962385, -1.4894602, 1.8407125, -2.9339611, -1.2927874, -0.7137091, 2.8515894, 0.6109025, 2.4848554, 1.1488599, 0.3455680, 2.1473437, 1.7231521, 2.1889389, 0.0262490, 1.6486843, -0.2450256, 2.2900939, -2.5290759, 1.9389485, 1.6840766, -2.3258119, 1.0110430, 2.6346169, -1.0978756, 0.1058508, -1.4360518, -0.2907172, -1.1895455, 1.0481918, 1.0516486, -2.0986858, -1.7708037, 0.7181241, 1.3296544, -1.3895290, -2.9396479, -0.8803832, -0.0595123, -0.2681628, -1.2932567, 2.8262648, 2.3084787, 0.9898864, 1.2336291, -2.3652806, -1.5707198, 2.7795698, -1.9976219, 2.9069782, 2.1887658, 2.8114732, -0.0850978, -0.3808674, -2.4582174, -2.9132564, -2.4653612, -2.1104009, -2.1344287, 0.6205779, -2.1846907, 2.2490064, 2.0779289, -0.2661282, 1.3820683, 1.6606495, 2.5595733, -2.0093659, 1.7549199, 2.1069071, -1.8321950, 1.3373799, 0.3379523, 0.7656077, -2.6763815, 2.1210568, 1.3261080, -1.0449514, 0.3755385, 2.4116810, 1.5713714, 2.6097816, -2.5386590, -1.8278706, 2.4162592, -1.0183215, -0.2284481, 2.8499867, -2.4355158, -0.0665855, 1.3785199, -2.3097419, -0.3298548, 0.7244548, 1.0877830, -0.2949900, 0.2998961, 1.5878361, 0.2986669, 0.4735249, 0.6635454, 0.9148462, 0.2126279, 0.3624573, -0.7084419, 1.4616585, 1.0493689, 2.9639192, 1.0662258, -2.0622934, 0.5767330, 0.0436070, -2.0912510, 1.8939626, -0.9901632, -0.8859261, -1.1236182, -2.3048336, -1.9347286, 1.0589359, 0.0824605, -1.8265792, 0.7583449, 1.0068165, 0.3427836, 1.3911102, 2.9031742, 0.7054775, 2.0568018, 1.3305605, 2.7597706, 0.7035823, 2.4407872, -1.5832443, 1.6857442, 2.3988490, -0.3984121, 2.8684415, -0.0522985, 0.0457977, -2.8228160, 1.4360643, -1.2429019, -0.2219502, 2.3959848, 2.6534356, 0.1432381, -0.6061285, 0.1442220, -0.8065366, 0.4853469, -1.3935527, 1.1326637, 1.1726874, -0.6500926, 1.4486285, 2.7468044, -0.4277649, 2.2339300, 1.9321610, -1.0290808, 0.4107683, 1.1324368, 1.6737951, -2.4523194, -1.9582967, -2.6961507, -0.2529235, -0.7776102, 0.3996878, 0.9231562, 1.3476469, -2.3787583, -0.9546120, 0.1145820, 1.5757079, -1.5889559, -2.8040414, 0.7327182, -0.5217076, 0.5566750, -2.2731884, -1.9974313, 0.2755160, 0.5696067, -2.1365977, -0.3532254, -2.6474783, 2.7128718, 0.2672850, -0.9057830, 0.4081128, 1.5191810, -0.8257630, 0.4799831, -2.2654271, 0.2700053, -1.5537992, -1.5798092, -2.4126486, 2.0430715, -1.3805383, -2.8643564, -0.5033156, 0.4146415, -0.1412935, -1.7395335, -2.7978750, 2.1043560, -2.4800572, 1.3317486, -2.4074284, -0.2518710, 0.6350209, -1.1808634, -0.5578050, -1.8559130, -2.0583397, 0.6041219, -1.1165436, 0.6863726, -1.1042814, -2.4586686, 0.6853267, 0.6004966, 1.9737566, -0.7577229, -2.9645475, 1.2513961, -1.0430615, -1.6968879, 1.2781859, 2.3237690, -1.5128401, 0.7459207, -0.3435556, -2.2745322, 2.1449100, 1.5411528, 2.9406002, 2.1085656, 0.0807730, 2.9226532, -0.6466167, -1.5559747, -2.7627878, -2.9430478, -2.7291211, -2.5928055, -2.8601551, 2.4387984, -2.3627559, -0.0150503, -2.6102146, 0.8649781, 1.0643224, -1.5247029, -0.6182565, 1.2536314, 2.8662587, -0.0329247, 0.4750775, -0.9715387, -1.9035549, -1.0914964, -1.3544170, 0.1828226, 0.1895280, 1.6646387, -2.2464576, 2.5008826, 1.8948309, -0.3062550, -1.5636466, -2.4023721, 2.5922414, -1.0565461, 2.3644604, -2.9229228, 2.8812776, 1.1622134, -0.7853366, -0.5243477, 1.4788846, -2.7662948, 0.7856511, 0.8022011, -1.5454869, -2.7528358, -0.8237265, 2.5237616, 0.1811504, -1.0015205, -2.0195119, -2.8408237, 2.4302389, -2.9259125, -2.0780823, 0.4890029, -0.6926393, 2.1168560, 0.9053710, 0.4579691, -0.8391535, -0.8394691, -2.5512823, 2.6008688, 1.4454133, 0.9034719, 1.2432188, -1.9347435, -0.2620923, -0.0521486, 1.0670932, -2.0212584, 1.5042146, 2.8825212, -2.5874754, -0.0868013, 0.1458466, -0.4638785, 0.1824468, 2.2324725, 2.8267777, 0.3899843, 1.7586414, 2.9471171, -2.3235328, 1.3577670, 2.5570990, 1.3327783, -0.4983757, 0.8434532, 2.3486153, 0.6140033, -1.5714422, 0.0013679, 1.3743619, 1.7742102, 0.9289980, -0.2992626, -1.7421640, 0.6195198, -2.5578436, -0.2576470, 2.8972402, 2.4323311, -2.5277921, -1.6135718, -1.1024422, -1.1958231, -2.6149399, -1.7180287, 2.9404201, 1.8097695, 1.1139174, -1.4919572, 1.7280718, 0.3186554, -2.2520714, 0.5191410, 1.7865163, 0.5591755, -0.5031777, 1.2325770, 1.8777689, -2.3950485, -1.5923735, 2.1303856, -0.1369453, 0.8089135, 0.7451434, 1.9434058, -0.5774685, 2.9667211, 1.3586573, 2.0442527, 1.9837300, 2.1751190, 0.4110373, -2.2615226, 1.5307801, 1.8930019, 0.3929919, 1.5971321, 0.6390496, -1.2351193, -1.0930796, 1.5854893, 0.9734172, -2.8040605, -0.0335031, -2.8195636, 2.1401887, -0.1024530, 0.2340937, 1.1451548, -2.2314893, 2.6731386, -0.1381867, -0.9054213, -1.3750292, 0.5243659, -2.4012682, 0.0398494, -2.5104690, -1.8016279, -2.4325307, -2.6224712, 0.8948087, -0.9491303, -0.9652882, -1.3860627, -1.1850943, -0.6410929, -0.8215726, -0.6404770, 1.9494035, 2.9216167, -1.0610194, 2.6254254, 2.0187504, 1.5223472, 0.0929619, -1.9111132, 2.8509312, -0.5933237, -2.5764571, -2.8776810, 1.4016783, 1.9048510, 2.1182437, -1.4448802, 0.1775361, -1.0258140, -0.7624929, 2.9510710, 2.1021871, 1.2191854, -2.3955153, -0.4262161, 0.9677978, 0.6803557, -2.6608914, 1.5070352, 2.5638578, -0.4506259, -2.7258424, 1.0674326, -0.4422243, 1.3353907, -1.9686388, 0.1814536, 0.5320421, 0.0252773, 0.1356287, -1.3820402, -1.0459860, -0.6307383, 1.7311081, 2.8257093, -0.0368254, -1.2298617, -2.4372063, 0.0355765, -0.8647202, 0.5190871, 2.9209275, -0.0920919, -1.2964846, 0.9085937, 0.6508892, 0.7693089, 1.3743779, -2.1079410, -1.7819069, 2.7178608, 1.2809284, 0.1521939, -1.5713562, -2.2621806, -2.8124930, -2.7123686, 1.7968505, 0.2740007, 0.7326887, 2.8967071, 0.6269129, -2.3016936, -1.7681540, -1.7989514, -0.9878778, 1.4327201, -1.6992400, 0.5979194, 0.6770967, 2.4864371, 0.3863588, 1.7642744, 2.8344400, 0.6901811, 0.4731531, 2.7016560, 0.2766846, 0.6407091, 0.6518424, -2.7558841, 0.1111460, 1.9772421, 1.1925030, -0.6214900, -2.2209254, 0.4157086, 2.9852318, -1.0791181, 2.0332461, -1.4889566, -0.6554831, -0.8112907, -1.9225915, -2.6955251, 1.4460746, -0.1321906, -0.8178164, -2.1512751, -0.8712213, 0.3957595, -1.6896418, 2.3245447, 0.5328237, -1.7690974, 2.6731490, -2.5190507, -1.3764308, 1.8379688, 2.3869520, 2.3291035, 2.2356117, -0.9046931, 0.8531967, 0.1547838, 1.3149609, -1.7495622, -2.1908248, -0.7237713, 2.4190304, -2.0734971, -0.3930996, 1.4507049, -0.5246662, -2.6504592, 2.9211344, -0.3073096, 1.7452790, 2.7204716, -2.9030686, -1.0564517, 1.4492554, 0.8740741, 1.8862460, -1.9254521, 0.7821477, -2.5615577, 1.5970232, -1.4967949, 2.4492791, 1.1157487, -1.6359090, -0.7777268, 1.7505647, 2.3110309, -2.1444463, -0.4129660, 2.0965677, 1.5914963, -1.6409403, -0.1286625, 1.4410403, 1.7598659, -1.8524580, 1.5203086, -0.3937422, 1.9902287, 0.2103905, 1.7262321, 1.6593291, 1.0296815, 2.2944848, -1.0480073, 0.8079307, 2.2305515, -0.6904688, -0.7389660, -1.8001770, 1.3218557, 2.8849964, 0.2137740, 2.4995356, 0.9949861, -2.8027641, 1.7593830, 0.3938029, -2.3627962, -0.6525126, -0.9791776, 1.3977479, -2.6361334, 0.0417210, 2.9007849, -0.1489020, 1.4909923, -1.9166968, 0.1100232, -1.8480977, 0.4300340, -2.7198915, -2.8565281, 1.9940950, -0.7715864, -0.1933993, -2.0098739, -0.3648774, -2.1798732, 2.0880526, -1.2375254, -0.6674027, -0.5597817, -1.1151654, 0.0442131, -1.9749833, 0.5064607, -1.5862074, 2.0985628, 1.1322721, -1.5146734, 0.4335653, -1.5237759, 0.8149226, -0.1192293, 0.0119451, -0.7802416, -1.9342581, -1.6826122, 1.7100933, -1.4751250, 1.2605082, 2.5212677, 1.7484698, -2.4782825, -0.4887095, 0.5315397, 0.8328367, 2.8556266, -1.5432819, 2.5682582, 0.4571400, 2.6862669, -0.5802469, -2.6939364, -1.1086469, 2.3455218, 1.5469815, -2.2422056, -1.7733159, 2.9971136, -0.8522183, 2.5013930, 0.1197851, 1.1834830, -0.5734159, 2.1919836, 2.6419044, 1.6987173, 1.7592407, -1.2878501, 1.8183318, 0.3744655, 0.5018163, 2.9970960, -2.8899352, 2.1591742, -2.0245610, 0.8976706, -2.4133824, -2.2449075, -1.2671278, 2.7791086, -0.6633154, -1.2647190, -0.8738263, 1.1496979, -1.5013543, -0.7438743, 1.6141336, 1.8280280, 0.8067328, 1.8503347, 0.9605673, 2.6742182, -0.1326146, -0.2562617, 1.7692080, -2.0276030, 0.5379532, -0.2354974, 2.7680389, 2.9511802, -1.9555834, 1.8972410, -2.9501441, 2.1434921, 0.7541654, 2.5012269, -1.8638570, -2.9814023, -0.3068554, 1.6653445, 2.7314312, -2.8142622, 2.4102096, 0.8809852, -0.4654641, 1.4563496, 2.9434186, -1.4999003, -0.1743871, 1.0524195, 2.9650689, 1.5651961, -0.6301778, 2.2280743, 0.7966274, 1.9367801, -1.5400866, 2.0777073, 2.6813166, -2.0077294, 1.5375985, -1.2967889, 1.4457946, -0.0469580, -0.8214340, 0.5976766, 0.9824620, 1.1886720, -1.5944337, -0.0752395, -2.4026915, -0.8017361, -2.8127794, -0.9895110, 1.0374106, 2.2179131, -1.3430752, 1.1321914, 0.5090396, -0.4671933, 2.1755665, -2.7295178, 0.6136583, -0.9364318, 0.6170572, -0.6723376, -1.2401303, -1.9953217, 0.6068312, -2.9824251, 2.9060533, 2.7291915, 1.2185972, -1.5226034, 2.2967394, -0.2902311, 2.3534816, -1.7682724, 1.6002640, -0.8782881, -1.3677393, 0.7020424, -2.3663983, 1.8948800, 0.1254733, 2.5983918, 1.3501658, -2.6953873, -1.9097422, 1.8830605, 0.5854587, 2.7160664, 2.5027222, -2.0921495, -0.4894772, -2.8422646, 1.8467036, 2.4560195, 0.2012036, -0.8646980, -2.3544088, -2.3125298, 1.6643058, -2.4835389, -2.8523854, 0.8022091, -0.1044182, 1.2696953, 2.4908175, -0.3920386, -0.8276511, 2.9621928, 2.1400584, 0.5549952, 1.2377685, -1.9612448, -2.4111212, 0.6909720, -2.5685791, 0.9709630, -2.6796797, 2.2588392, -2.1684219, -0.6444365, -0.1215344, 2.3563169, -0.5577174, 0.1909969, 0.1478876, -1.7038561, -1.7651639, -1.0461539, -1.7861204, -0.1391173, 1.3595511, -2.6738626, -2.7083848, -0.3810618, 1.0479041, -2.9750720, 1.2961766, -0.3018671, 0.0893071, -2.7213102, 0.3258295, -2.7113712, -1.1566498, -0.3027197, 0.3388289, 2.4379423, 2.2255459, -0.3270102, 0.6981937, -1.7066905, 1.5311677, -0.9807049, -1.9590964, -2.4075168, 1.1166960, -1.8583796, -2.1426665, 2.2010506, 1.0494119, 2.7483607, 2.6410494, 0.4636387, -0.0294706, -2.9342550, 0.2548406, -2.7797663, 0.9649637, 1.3699188, 0.1353873, 2.4059810, -2.2859978, -1.7007175, 0.5687648, 2.3470417, -1.8459383, 2.6415981, -0.0552869, 2.2329112, 1.6942133, -0.0273283, 0.8787984, -2.8029297, -1.5270497, 2.6365407, -1.4387712, -2.5338779, 0.0077031, 2.6546550, -1.6363444, 0.7004331, -0.8109421, 2.0195242, -2.4256822, 1.2325685, -2.8438105, -2.6108863, -2.4443646, -2.2798197, -1.2159075, -0.4257529, 0.4565495, -1.4599001, -2.5236877, -1.7226515, -1.3408532, 1.5679127, 1.4960705, -1.1976537, 0.9647072, -2.2341619, 0.6281540, 2.3425684, 0.6707865, 1.0489656, 0.4033546, 0.4764383, -1.7657270, 1.0028224, -0.3849607, -2.0991703, 1.3097452, 0.2286620, 0.9864063, 0.7246606, 1.0289193, -0.2946667, -0.0724575, -2.2199466, 0.4177591, 2.6847237, -1.4113425, -0.3161552, -0.0703902, 0.2270945, 2.3326625, 2.7325843, -1.8579023, 1.5854183, 2.0869367, -2.7069394, 1.7998324, 2.2658385, 0.4676389, 1.3642862, -2.2087792, -1.0047102, 2.6688860, 1.9703556, -1.2398487, 0.5052389, 2.7645168, -0.1001429, 2.8286802, 0.7168955, -2.5411502, -2.5866323, 0.7145215, 2.2886295, 1.0951219, 2.3009466, -1.5982364, -0.6333588, -1.6944915, 0.0861095, 2.8005112, -1.3034459, -0.3232764, 0.7338714, 2.8328320, -2.1368351, 1.8600435, -1.8539840, -0.0230579, -1.6318515, 0.0996541, 0.9862747, 0.0419532, -0.5346216, -2.3873002, 0.3321532, -1.2106828, 1.1171760, -2.1181312, 1.8657160, -2.3131628, -2.1818099, 2.8766598, 1.7197253, -2.2186212, -2.9860425, 2.5181754, -0.0361523, -1.7636521, 1.1003684, 1.4390359, -0.0566613, -2.8198700, -2.3655885, 2.2902953, 1.8875163, -2.5572968, -1.3318183, -0.4094399, -1.0210498, 1.7273730, -2.1331164, -2.7770935, -1.3223928, 0.6811583, -2.7458085, 0.3161231, 1.8016334, 0.9914056, -2.4622687, -2.3827795, 2.2666485, 2.1846297, 1.5066912, -1.4201912, -2.2975734, -1.5628956, -2.7408895, -1.9982376, -1.1891011, 2.2377457, 1.0181842, -1.0897571, -2.1034054, -2.4482188, 2.5056895, 0.3511995, -1.8392622, -0.9828376, 0.8136923, 2.8453706, 1.3778958, 2.8601277, 0.5258072, 0.9247059, -0.7731391, -1.3063799, -2.9727249, -0.6816919, -0.5084319, -2.1322878, 1.9210401, 0.4276066, -0.3886493, -1.6833672, 1.3908485, -2.5433985, -2.7468386, -1.2111254, -1.6207504, 1.5087053, -1.2777977, -1.6640738, -2.3638791, -0.5767014, 2.0828081, 1.2003268, 0.7436836, -2.5065555, -1.1740368, 1.5201164, 1.4409965, -2.9861396, -1.8301814, 2.8516659, -0.1597438, -2.2658427, 2.1154637, -1.2640472, 1.7967612, 2.8556653, 0.3493088, -1.9729704, 0.8172176, -2.4091823, -0.3949451, -1.4644254, -1.6940051, -2.8879392, -2.4396984, -1.9410484, -0.7070812, 0.8450399, -0.2692975, 1.8269176, 2.7589627, -2.5092032, 2.1695690, 2.1551012, 2.2849190, -0.7361100, 2.4704795, -2.2696875, 0.6213761, 2.8716662, 0.4229031, 1.3680266, -0.0510994, -2.3114240, -1.3578101, 2.4586691, 0.1157782, 1.1689915, 2.0804137, 2.4180088, -0.1565325, 1.5085152, 1.4875653, -0.2651245, -1.9627576, -1.7843571, 1.7419973, 2.1782114, -1.5256899, 0.4979692, -1.1170096, -0.1259374, -2.0871751, -0.9345161, -0.7792924, -0.0338203, 0.7602205, -0.7081150, -1.4680059, -1.1950200, 2.2663775, -1.1399934, 2.3554419, -1.1943484, -0.7671867, 2.1130748, -0.7291957, 2.9846901, -1.7589413, -0.1571630, 2.5286697, 1.4943674, -2.1902516, 1.6840268, -0.4795781, 1.6920219, 1.8094572, 1.0084843, 1.9193450, 2.0950883, -1.3450089, 1.8504568, 0.6943711, 0.7515080, 1.3527875, 2.1786956, 1.3684516, 1.7680779, -0.1750171, 2.5377590, -1.2700084, -2.3509088, 0.6067816, -0.6830878, 2.8527470, 2.5612720, -2.4957681, -0.8539531, -1.5945497, 1.9274479, 1.7547248, -0.1402884, 2.9601131, 0.2663657, -1.5480808, -2.1055150, -2.9259754, -0.4918357, -0.2821437, 0.5853145, -1.2386257, -2.6513605, -2.1983273, 2.3430038, 2.9619328, 1.0689081, 1.7337883, -0.4614221, 2.6865920, 0.5568551, 0.2753873, -2.0575216, -1.7141308, -1.0743417, -1.7045182, -0.6176617, -0.8644747, 0.0989876, 2.6536880, -0.8901545, -0.5791442, -2.2777106, -1.2473826, -2.1557455, 2.7239186, 1.8004861, -2.8418633, 0.7296647, 1.6565949, -2.9699832, 2.0717528, -0.8740516, 0.6695554, -2.4356069, 0.5028589, -0.8579409, -0.6766667, -2.0709091, -1.6806184, -0.1174674, 0.6037802, 2.3693628, 1.9737036, -0.4760657, 2.5686586, -1.8651941, 0.4818700, -0.7715486, 2.2211621, 2.8785342, -2.8458088, 0.6124073, -2.6139795, -1.3179420, -2.2029176, 0.7122504, -0.6372066, 1.7047626, 0.2947832, 2.2381895, -2.3870256, 1.5279716, 0.8950577, -0.8656229, -1.0121953, 1.6480785, 2.6960101, 2.5832098, 1.2649772, -2.6429419, -2.6369479, 2.4439179, -2.1311944, -1.8649726, 0.5170970, 2.1734756, 1.1859563, -1.4256789, 1.4206125, 1.5395699, 2.3417582, 1.1011784, 2.9765894, 2.6883504, -2.2831685, 2.6022868, -0.5784911, -1.3332894, -1.7339985, 2.3865027, 0.5877928, -0.5259110, 2.4610879, -0.7384727, -2.0247247, -2.9498303, -2.0878667, -2.9279557, 0.2205644, -0.6319052, 2.6301226, 0.3628394, -1.0635184, 2.1977212, 2.9401780, -1.1486708, 1.8499575, 2.6947895, 1.3953492, -1.7965508, -0.1383138, -0.9429915, 1.8362512, -1.2636350, -1.5095135, -2.2488659, -2.6588723, 2.7496549, 1.8456856, -2.6596136, 2.4782517, -0.3907147, 1.6706669, 2.4387148, -0.8014566, 2.8261752, -0.6908051, 0.2160163, -0.6580837, -0.9893022, -0.2466997, 0.2870313, -1.2009623, -0.0617822, 0.0514868, 2.3984757, 1.9784981, 2.6646227, -1.2669396, 1.9780462, 1.3112294, 0.0829331, 2.7375250, -1.9311317, 2.6047991, 0.2509232, -0.5442298, -2.7914033, 0.0957567, -0.5715891, -1.4431296, -2.0687319, 1.3946545, 2.1301337, 1.8106224, 1.9612128, 0.9768127, -1.8650752, 2.5621034, -0.7054044, -0.2982698, 1.4220184, -0.7981440, 2.2125742, -1.3550281, -0.6150118, 2.5240198, 0.5351237, 1.9901329, 1.5182435, 0.7622156, 1.1086326, 0.2689197, 2.0547433, 0.2355680, 2.2179909, 2.0052606, 0.3402738, 1.4952713, -1.2343806, 1.7990392, -2.1919852, 0.2948511, -2.5522444, -2.7838811, -2.7385508, 0.8215394, 1.4816778, 1.2864857, 0.8512044, -1.9381330, 1.1203740, -1.2954545, 1.2013250, -1.3379309, -1.1931150, 0.6136999, -2.2461464, 2.5192240, 1.4226769, -2.1164976, 0.3126372, 1.0568031, -2.6176638, 1.0369280, 0.7884688, 2.6079790, -1.4036015, -0.5045465, 2.5258302, 2.4089685, 2.7963947, -0.8598630, 2.4019716, -1.5955648, 1.3362458, 0.7976548, -0.4821074, -1.7171970, -1.6140491, -1.2869797, -0.8303064, -1.7455844, -1.7339812, 1.7989021, -1.8656641, 1.2476984, -2.5118471, -2.8852696, 1.8637037, 0.8787365, 2.4229245, 2.4993289, 1.7914183, -0.7298639, -2.5504608, 2.4692817, -2.8066371, -1.9982474, -0.7521202, -0.8502294, 1.8655134, 0.5705702, 1.6033495, -2.6361846, 2.0733974, -0.7406194, -1.3451911, 2.9977786, 0.1742250, -2.3649225, 1.2638071, -2.7343437, -2.8950113, -2.2533654, 1.4453294, -2.1756806, -2.0918913, -2.3507059, 1.4535570, 2.3970910, 2.6101861, -0.0593780, -2.7243139, -1.0296179, -0.8180302, 1.9479053, 0.6400131, -1.7844643, 2.1444027, 0.2316566, 0.1798395, 2.6890468, 0.1803159, -1.6218768, -1.0142068, -0.4611843, 0.7974169, 1.6437731, 2.7363038, 1.7578842, 2.4564751, 0.9308821, -2.4097756, 0.0820701, -0.5599522, -2.7775390, -2.7901535, 2.2673857, -2.9995990, -2.6004645, -0.3867230, -0.9017631, 0.4622522, 2.3497809, -2.4286312, -1.7033386, 0.3415659, 1.8968897, -1.1155816, -0.1251515, 1.7794046, 0.7669365, 0.5887400, -0.8642081, 0.4835992, 1.1487305, 2.7891299, -2.0170869, 1.6167429, -2.0567841, 1.6340642, 0.3108321, -0.1472037, -2.5267298, 2.6365190, 0.9529433, 0.1161744, -2.9175805, -0.7114283, 0.1155190, -1.8569342, -2.3798481, -0.9368807, -0.7176997, 1.6131455, -2.5353141, 0.5816953, 1.8928584, 1.5017115, 2.8125911, 0.1312774, 2.5472660, -2.3110951, 0.9388813, -1.2940127, 1.1650295, 2.5903607, -1.5773351, -1.7772706, -2.7340188, 2.6782573, -2.3625498, -2.4034447, -1.1201185, -1.9250056, -0.6679811, 2.4158735, 2.6761730, -2.5132234, -1.4786331, -0.8463218, -2.1479285, -1.1705251, 0.0850684, 2.0419293, -1.7076416, -0.6817852, -1.2606182, -0.5921929, -1.0257683, -1.0036710, -1.1125311, -1.4009623, 0.7706870, 0.1920046, -1.2970770, 2.7743931, -1.5399109, -0.2942965, 2.6145593, -0.1377926, 2.8645804, -0.5069271, -2.4551715, 2.5533144, -2.8729503, 1.6897709, -1.5593906, -1.2336522, -2.1699377, 0.8371981, 0.5539656, 0.0491114, 0.6413405, -2.0331800, 0.5191277, 2.6204472, -2.7225191, -0.7408618, -0.5962089, -0.7057325, -0.3653331, 2.1434452, -1.6240164, -2.7507732, 1.0324172, 1.3209125, 1.0850150, 1.4115223, -0.3477202, 0.9460749, 2.8210246, -2.0035021, -2.7405420, -1.9493204, 1.3227381, 2.1625560, -0.7689359, -0.9813059, -1.2134851, 2.2341451, -2.4233665, -0.0308664, -1.6829601, 2.3141064, -1.3080537, -0.5991352, 1.6581045, 0.1512865, -1.8015222, 2.7822114, 1.1434465, -0.5297533, -0.1647487, 0.0866091, -1.1915943, -2.7943459, -1.8131111, -1.1273486, 0.1566885, 1.6977738, 1.6688928, 2.2294954, 2.7279748, 0.2412541, 0.7348725, -2.7351347, 2.3070445, 0.1288354, -1.2759624, 2.8447572, -0.3994257, 1.0685497, -1.3569444, -1.8400874, -0.3538517, -1.5564054, 2.0738164, 0.0525100, -2.7696363, 1.5057201, -2.4752244, 0.9412938, 1.4423158, -2.0601549, -2.8933591, 2.2958444, -2.7571537, 2.1849178, 2.5413152, 2.8721506, -1.0155003, -1.7722072, -1.7214847, -1.8629140, 0.2138528, 2.2087543, 0.5999905, 2.2216390, -2.6495484, -0.2868093, 2.8973666, -0.6660620, -1.1196735, -0.1582930, 0.3684290, -0.3437574, 1.9117714, -1.2888665, -0.7514117, -0.5333452, 2.5415053, 0.3275731, 0.1454252, -1.5599920, 2.1640988, -0.5862613, -1.8195464, -0.9662896, -1.3160864, 0.2248350, 1.8205341, 1.9164644, 0.8961342, -0.5295498, 1.9842921, 2.8817919, -0.8478583, -0.5717988, 1.0155429, 0.6659084, -1.8910657, 0.9459179, -0.7516965, 1.0808439, 2.1776376, -0.7245122, -0.3642357, 0.1475644, 2.7297274, -2.1247870, 1.1625888, -1.8112999, -2.2234060, -1.2116120, -1.5064390, 0.2742734, -0.1874601, 1.4041202, -1.9495366, 2.0627301, -0.6856274, 2.2086845, -1.6854089, -0.5036245, -1.0066884, 0.1487738, -0.4752217, -2.5922061, -0.9735073, 2.7229877, -2.2199356, 0.5665673, 1.5473607, -2.4901120, 0.1658889, -0.6220414, 0.2693217, -1.2406119, 2.6040253, 2.4381387, 2.2942447, -1.6948012, -0.2475712, 2.2267201, -0.6997538, -1.7270588, -2.3573673, -1.8600510, 0.9663675, -0.1266671, -2.0543145, 1.3075002, -1.5475751, -0.5324963, -0.8764474, -2.6528207, -0.8233309, 0.1071103, -1.6216904, -0.8596169, -1.2679241, 0.5832066, -2.7515183, -2.9122922, -1.1661014, -0.6843847, 2.7971512, 0.5006971, -1.3112215, -0.4154407, -2.4635666, 2.7552851, -1.2706375, 0.5202134, -1.3961929, 1.3269307, -1.8290414, -2.6043199, 0.9725119, -1.8262118, -2.2105422, -2.0807926, 1.1893274, -0.9334613, 0.3493687, 0.5992853, 1.3611848, 0.7083457, -2.0769094, 0.9976851, 0.5370498, 0.4040142, 1.2941336, -2.9241476, 2.5946371, 2.4773858, -2.2023106, -2.6384661, 2.8614238, 0.4025413, 2.9183363, 0.8159053, -1.8104248, -1.8149928, 2.6478337, -0.9438817, 2.6751722, 0.2419408, 2.2821225, -0.0023988, -1.2743947, 0.9663042, -2.9199260, -1.4833955, 1.6156723, 0.5354713, 0.1346021, -0.4110949, 0.6310810, 2.1095885, -0.3341059, 2.3658160, -2.7691844, 1.3349417, -2.5590342, 0.0048543, 1.4103619, -2.7639982, -1.8754867, 2.1625426, 0.2657096, -1.4067256, -1.6703469, 1.4222083, 1.6468911, 1.3092465, -2.6684191, -2.8043254, 1.6809303, 1.2792164, -1.6341245, 0.2756793, 1.4003428, -0.3555607, -0.1795459, 0.8925883, 0.9475000, -1.5446242, 2.5260674, -0.4922688, -1.0615911, 2.8899053, -2.5756429, -0.7282354, 1.8372147, 0.6035019, -1.3847911, 0.4137018, 2.2192853, 0.4652544, 2.8147264, 2.7135985, -2.1700565, -0.2654118, 0.6841956, -1.4167603, 0.5185653, 1.9990160, 2.7159680, 0.6106689, -0.9394354, 0.0802520, 2.8876278, 0.3563469, -0.2006326, -1.7295009, 0.3609733, -0.5068000, -2.1428475, 2.1948683, 2.0317037, 0.0821128, 2.3190338, 1.0178069, 1.0415177, -2.2063970, -2.7186830, 0.5717487, 2.2099332, -2.5548259, 2.2144717, -0.9450383, -2.7210332, 1.3594545, -0.0887004, 2.6186503, 2.0998987, 0.8048175, 2.3951136, 1.6980036, 1.6678999, -1.4210785, -1.9202056, -1.6613541, 1.9659724, -0.0470127, 1.2272544, -0.8810207, -2.2892635, 2.2688047, 2.6622784, -1.4058050, -0.8244499, 1.9050493, 0.1488014, -2.8737789, -2.1608657, -2.6809973, 0.2483631, 1.3828571, -1.6468005, 0.6916970, 1.7750776, -1.1256782, -1.7734390, 2.4303634, 0.4060812, 0.7255712, -2.2153918, -1.0425311, -1.2881107, -1.4613270, 2.0664224, 0.5566274, -0.3627693, 1.2546990, 1.6851310, -0.0988651, 2.2138602, -2.1696786, 2.9310572, 1.0789740, -2.9217237, 1.9331874, -2.0491083, 0.3839593, -0.8117780, 2.9962094, 0.2543000, -1.2145919, -1.3026483, 0.4859838, -0.2526482, 1.8628376, 1.2505691, 2.7711923, 0.4744236, 2.4924172, -0.9423320, 0.9269377, -1.7015076, 1.5920308, -1.8435930, -1.6971753, 1.0554321, 0.5263756, 1.5965719, 1.5783155, 0.8781420, -1.6523942, -1.2164452, 0.8115856, 2.1160490, 0.0007448, -2.9058001, 1.6419030, -1.9168740, 1.3007380, 1.7557200, 2.8455186, -0.3044893, 1.7267452, -2.4279685, -0.0919103, 2.3841604, -1.4779264, -0.2526709, -2.9969114, -2.6205681, 2.0169124, -2.8422437, -1.3567874, -0.5377871, 2.5881821, -2.1308124, -2.2779771, -0.3432010, -1.5678719, -1.9905287, -1.5188148, -1.4894789, 0.1007286, -0.9767712, -0.0669824, -0.0446031, 1.6409563, 1.4364323, 1.0465701, 1.7982306, 2.8562486, 0.2955264, -0.2066594, -1.4944161, 0.5551314, 0.8923335, 0.2694081, -1.4294558, -2.0516577, -0.7086111, -2.6847841, -2.3295590, 2.3957610, -1.7305361, -2.8395329, 2.3316958, 1.1303728, -0.2269145, 1.8661900, 0.4579452, -1.2890298, 2.3053829, -1.3077782, -2.4297114, -0.2624895, 2.1100661, 0.3453218, 1.8066004, -0.8387052, -0.3235317, 0.0223006, -2.2402402, 1.4198936, -2.0841971, 0.1770885, 0.4883532, 2.8219481, 1.6357015, -1.2988670, 2.8637593, -1.8387818, -2.4298745, -1.9788106, -0.7059397, 1.4850229, -1.9427012, 0.3980459, 2.3436530, 0.7246171, -2.6383597, -1.7264796, -0.8144007, -2.6236401, -0.4477839, -0.7837906, 2.4947082, -2.1507623, -1.5455607, -0.5308454, 1.2613268, 0.4010762, 1.3637586, 2.6240603, 1.9873096, -2.5055930, -1.9406688, 1.0547723, 0.5320650, -1.3327140, -2.4719083, -1.2710623, 2.3543169, -1.7342992, -2.8695921, 0.3352985, 0.1584703, -2.7424820, 2.1511685, -2.1343076, 2.2202792, -0.4329429, 1.5733276, -1.9719279, -0.9399342, -2.0931870, 1.6898283, -0.0021654, 0.3147535, 1.1770285, 2.0749488, 2.8738905, 2.1681918, 0.6605337, 0.4020113, -1.1128598, 0.4277010, -1.1562678, -2.5103723, 1.0947359, -1.1155828, -2.8766537, 2.9921036, -0.0506574, 2.8182073, 0.0315965, 0.3724173, -2.9878129, -0.8608847, 0.6159394, -1.2844526, -1.3516570, 1.2558639, -2.0209142, -2.2746110, -2.6017259, -2.7877740, -0.5806906, 1.5506008, 2.3493073, -2.8097797, -1.4798654, 2.7544720, 1.2061076, 0.6062914, 0.7631951, -0.0032604, -1.4381828, 1.2740515, 1.9373495, -0.2688742, 0.6619865, 2.8362266, -2.4464909, 2.6892525, 0.7922363, 1.9314759, 2.7616387, -1.9535308, -2.8291724, 0.4389820, 0.0293761, 1.2227168, 1.1894766, -2.5814198, -2.2323565, 2.8098710, 1.1292484, -2.5397510, 1.4026213, 0.1074786, -0.6209388, 1.5380973, -0.1127171, 1.5689853, 0.1825242, -0.1906479, -0.2429834, 1.7849657, 0.4846407, 2.1783367, 1.5674416, -1.0911242, 1.6036358, 0.2483815, 1.7317833, -1.0357052, -1.4058814, -1.3128256, 0.5917013, -0.1731844, -2.3195791, -2.3747455, 2.1475663, -2.2732406, 0.4568391, 1.7830073, -0.7874368, 0.7798410, 2.5620837, -1.9511504, 0.6380295, -0.5942617, 1.2076578, -1.9983536, -1.9786035, 0.9888323, 1.5633405, -2.9737529, -2.6870661, 2.1354501, -1.8239319, -1.8628359, -2.5467091, -1.5989408, -1.0309129, -1.3061225, -1.1018318, 2.4394684, -1.9809355, 2.2969194, 0.5028592, -0.8934745, -0.4307358, -0.6911573, 2.0788407, -0.6435813, 0.4601009, -0.0362326, 0.3843259, -2.9083573, 0.4108905, -2.3033187, 0.5139394, 2.2406361, 0.2017796, -1.8351377, -2.4004009, 2.5287433, -2.6218114, -0.2250874, -1.9915447, -1.4398613, 1.6948779, 2.5515185, -1.8223085, 2.9695506, -1.8671375, 2.9543165, -1.4957068, 1.1504710, -0.2735792, 0.6699419, 1.5148182, -1.8912635, 2.5589411, -1.9977945, -0.0025640, -1.6144656, -1.5738929, -1.8495038, 0.3282155, -2.8306140, 0.1725178, 2.6445464, 2.6768158, -1.1846320, -1.5727172, -1.5313007, 0.8288604, -2.1500217, 0.6892216, -1.0334337, -2.5971550, -0.0223717, 1.5606428, -0.2908582, 2.3666334, 0.3335127, -2.9185962, 0.3382638, -0.6008942, -0.2681314, -1.8379904, -2.7645702, -1.1846706, 0.1777577, -1.8817107, -1.4187996, -0.0704601, 1.3578506, 1.7095701, -2.7984389, 0.7037300, 2.7836198, -0.6974443, 1.8482659, 1.3202456, 0.8557717, 1.0933333, 1.0809805, -1.8837371, -0.0046733, 0.8971151, 0.0423735, 0.4816638, -2.8543441, -0.7725330, 2.8788760, 2.4533293, 0.3663479, 1.6613392, 2.8359479, -0.8620768, -1.6410102, -0.4171476, -1.9405209, 1.0592961, 2.5392154, -1.9907719, -2.8840830, -0.3485550, 2.0009677, -0.0627835, -0.2606764, 2.0418762, -0.5052335, -1.3896663, 1.6297399, 0.4190859, 1.9472197, 1.0657707, 0.1526798, -1.4305537, 1.2097277, -0.5129570, -1.6593185, -0.4854500, 2.7999061, 0.2906135, 2.6991658, 0.5839462, 1.9805157, 2.6613285, 0.0008217, 0.5715020, 1.3624693, 2.1069151, -1.8301483, 0.7196101, 1.0187688, 1.9271943, -1.3176431, -2.6752592, -2.0482208, 0.4866627, 1.2888337, -0.6400002, -2.3304061, 0.7579826, -2.1979348, -1.6567940, -2.5113246, 0.0175368, 2.2588033, 0.6709822, -2.6445147, 2.7284858, 1.7171867, 1.0193756, -2.9702046, -1.7278458, -2.8871148, -1.7472779, 2.5087253, 0.1824202, -1.8942040, -2.4732474, 2.7284799, 1.1469567, 1.4230088, 1.3917025, 2.1919196, -1.0936275, -2.1442708, 2.7923223, 1.4596341, 0.3014173, -2.9303889, 1.0216058, 2.6525811, -1.2233484, 1.3045694, -1.2232799, -0.7886695, 1.5805408, 1.5529944, -1.0529403, 2.5509673, -0.9625454, -2.2556310, -1.1010229, 0.7113281, -1.5524885, 2.3288328, 0.4569275, -0.9936717, -0.4014956, 1.6800755, -2.6221955, -1.6664482, -2.3191911, 2.9068015, 0.2292843, 2.5263565, 0.2566813, 1.1108026, 1.4739815, -0.1107100, 1.6042402, -1.1589909, 0.8275380, 1.2560952, -2.9037793, 1.1817076, -2.3712832, 1.0073693, -2.1992404, 0.2332419, -0.5661812, 2.4333481, -0.3610500, 2.5573253, 1.7885675, 0.5659787, 2.0817053, -0.4243075, -2.7731803, 2.3313119, -2.5786895, 2.1633545, -1.1721687, -2.6005992, -2.8759871, 0.7134312, -2.5278291, -1.7295633, -0.9295371, -0.3636054, -1.9032781, 0.7262806, 2.0311773, 2.7243584, 0.3041706, -1.3561573, -0.8691931, -0.9944722, -0.3456383, -1.4212470, -1.6859234, 1.7744781, -1.6975574, 2.3383131, 2.9438775, -1.9664829, 0.4393397, 1.4237842, -0.1976952, -0.2840862, 2.0621616, -0.4939772, -2.7985402, -1.4092642, 2.8407849, -0.5403961, 0.5739071, 1.6438624, -1.5242112, -0.5423296, 2.0504805, -0.3911678, -1.9900540, 1.8904825, -1.4584982, 0.0300343, 2.3499946, 0.4000232, -0.7554957, -2.3882501, 1.1892251, -0.6129164, -2.9182853, 1.3035287, 1.8782252, -0.6656963, -1.2744550, 1.8792085, -1.2704281, 1.3417571, -1.4677357, 1.0723585, 2.1540617, 0.0514082, 0.7136867, -2.4740674, 1.2546301, -2.9685725, 1.5744123, 0.6274219, -0.8407106, -1.1670041, 2.5665319, -0.5447482, 2.0391592, 2.7021256, 2.2037865, -2.0604517, 1.4727257, 2.0891287, 1.4395275, 2.2171862, 0.0263808, -1.4362017, 2.3129550, 2.2532611, 1.2988049, -1.2154211, -0.7828437, 0.1681206, 0.3326136, -0.9495644, -2.3677403, 0.9219108, -1.0484028, 0.5466104, 2.8262220, 1.7944245, 0.9329804, -0.4122116, -1.3254542, -0.9192786, 0.0175422, 1.7424898, -2.4799929, -0.3578409, -0.6781863, -2.2103974, -2.3721424, -2.7226572, 0.2590171, 1.2129088, 2.0180181, -1.7052326, 0.7679690, -2.0021709, -2.5372597, -2.2406920, 2.4134854, 1.1585720, 1.5457010, -2.3122292, -1.3030695, -2.6131240, -1.5778555, 1.2500387, 2.6388644, 1.9216734, -2.0403661, -2.4527913, 1.1471990, 2.1108353, 1.6990254, -1.6612493, 0.1631717, -1.5654288, 2.4617087, 2.5060070, 1.6620362, 2.4731263, 2.8157617, -1.8706300, 0.7059425, 1.2232238, 2.6915280, -2.5822037, -0.6998616, -0.2085932, 0.7826689, -2.2644197, -1.5178664, 1.6650439, -2.8556517, 2.7809253, -2.7851610, 1.4279469, 2.4005334, 1.4138738, 0.9039012, -0.2964155, 0.1558428, -1.2648219, -1.1058231, 0.3191149, 2.1959812, 2.2617634, 2.4032604, -0.9738350, 1.6531128, 0.4560531, -1.5896441, -2.1624927, -0.6655449, -0.9388425, 1.7768405, 0.5632959, 1.7217865, -2.7055529, -0.6167032, -0.8330071, -1.1162942, 2.2295774, -1.3306736, -0.9426314, 1.5187503, 0.8400782, 0.3309263, 2.7745761, 1.1281283, 0.2992539, 1.3185562, 0.1023612, 2.8316911, 2.9670347, 1.8504271, 0.5892527, 1.5712330, -2.9158207, -2.8519611, 0.2685535, 0.7708400, 0.9099256, 0.9870705, 0.6454166, -2.7507849, -2.4922216, -2.0230717, 2.3935758, 2.6268277, -1.6823587, 1.3437759, -2.7733739, -0.8291315, 1.9217601, -0.5178864, 0.4349355, -2.2856629, -2.6631730, -0.1728816, -0.3552105, 2.5167691, 1.9167724, 2.0709802, 0.2045255, -0.5987474, -0.5025611, 1.2480488, -2.4046614, 2.7349633, -0.9620913, -0.0973747, 2.3770360, -2.8352273, -1.9903691, 2.3971832, 0.6549449, -0.7835920, 0.1501708, 2.8958347, -1.7711385, 0.7645424, -1.2121822, -1.9665348, -2.3432530, 2.3971652, -0.4328786, 2.4848856, -0.0376304, -2.2760751, 0.8146395, 0.2813588, 0.8561186, -1.4776160, 2.9564403, -1.5131028, 2.1964046, -2.2343066, -2.6199315, 2.2590939, 1.0978945, -1.7073014, 1.6307651, -1.0998716, 1.7641913, -2.7446649, -2.7894070, -1.7437922, -2.8761559, -0.8195690, -2.0855428, -1.2654415, -0.8756672, -0.6884301, 1.2219698, -2.1330904, -1.4014325, 2.7151633, 1.8485813, 0.9941381, -0.0573087, 0.2849044, -1.0249640, 0.9942162, 0.4263953, 2.2106300, -1.2485216, 2.3095773, 1.5642528, 0.8729572, -2.2630198, 1.7963833, -1.0785230, -1.7521439, 0.5563552, 0.6897372, 0.4537577, 1.9734736, 2.4283902, 1.6113801, 0.5719196, 2.1097589, -0.7375283, 2.9992164, 2.1608185, 2.9728138, 2.8096462, -0.6022524, -0.0393498, 1.0839911, 0.9983712, -2.6564259, 1.0075773, 2.1380520, 0.9952343, 2.1008520, 1.1729479, 2.6541938, 1.3418215, -2.1272846, -1.3105605, -0.4361264, 2.2249632, -0.7150609, -2.7825930, 0.2672931, 0.1567250, -0.3364321, 1.0362660, 2.3112379, -2.3847745, -2.1593520, 0.1856160, 2.5973286, 1.0472533, 1.0396870, 2.9566243, -2.0062837, 0.2913448, 2.7498115, -0.9488732, 2.6076517, 2.6533435, -0.8103888, -2.4410273, -2.9196372, -0.1517497, -1.1088591, -2.9964508, 2.5045781, 0.7569881, 1.4661998, -0.6525191, -2.9446412, 2.9202523, -1.6279579, -1.7439915, 2.5908097, 1.8706381, 0.6452040, -2.6312718, 0.5142970, 2.2628782, -1.9458449, -1.2974447, 1.4043532, 0.1980647, 1.9155800, 1.7266731, -1.9991198, 1.7540814, 1.7586237, 0.1134789, 0.2847834, -2.9699682, -2.7422511, -2.8903712, -0.7397238, -0.6028730, 1.8502944, -2.9230680, -0.3820375, -0.0170045, -0.8973363, 1.3218629, -0.8635567, 0.8402188, 0.1348298, -0.1221881, 2.5943097, 0.1412209, -2.2414827, -1.2364283, -2.7165304, -1.0634163, -0.3436664, -2.2269077, 1.1371890, -0.3858606, -1.5126306, 0.8723747, 2.6708711, -1.3082505, 1.5768930, 1.4363255, 0.8394500, 1.2432843, -2.9264464, 0.5786551, -1.0976110, -1.4595363, 2.5051444, 0.6708679, -0.9862948, -2.9433870, -0.9863415, 2.7488171, 0.9110892, -2.6745390, -2.2778992, -1.0182481, 2.7298934, 2.1296119, -2.6124427, 1.9438389, -0.2770393, -1.8535605, 2.7311726, 1.8179660, -0.6433435, -1.5311525, 1.4903827, -1.2664725, -1.0239257, 0.6392857, -0.4851807, 0.3274647, -0.1788449, 0.0031309, 2.5515423, 1.0146344, -2.8498779, -2.1816105, -2.6942156, -2.8155830, 2.8111383, 0.8154767, 2.4815386, -2.0004990, -2.6706870, -2.9093033, 1.3383483, -2.0404897, -1.4206539, -2.0979401, 1.7600641, -2.1329996, -1.8693565, 0.1643868, 1.9649430, -2.9118802, 2.6059558, -1.6941197, 0.0503791, 0.7117063, 2.9585682, 0.1035052, -0.5465091, 0.6296814, -0.9343340, 1.7130294, -2.9187675, 0.0813767, 0.0731775, 1.1031662, 2.6149603, -0.0377079, 0.8702296, -1.4599108, -0.8347059, 0.1039918, -0.1552329, 2.5813503, -0.8545132, -2.9688290, 2.7691915, 0.0669167, -2.2383567, -2.8225872, -2.9861204, 1.8115394, -0.3895370, 1.4619770, -1.2882640, -0.4366751, 2.8143602, -2.3931363, 1.7405013, 2.6510297, 1.9577557, -1.5021537, 1.0497642, 0.3622563, 1.3014565, 1.0976787, -0.3753163, -2.9673187, 2.4674228, 0.7654221, -2.6143071, -1.3001185, 2.4478609, 0.4781559, -1.0395563, 0.8498183, 1.5468708, 2.8410277, 0.7140691, 2.8192225, 0.6257489, 2.3561852, 2.2542674, -1.8531548, -1.7457163, -2.7326262, 0.7193246, -0.0767482, -0.4501014, 0.7147772, 1.9250761, 2.1149062, 1.8951221, -2.5336170, 1.9325083, 1.8133279, 1.5808182, 0.9762821, -2.8470950, 1.9412443, 2.7174785, -0.1327586, -1.1295681, 1.4994888, -1.4378618, -2.0711128, -0.8911860, 1.5914936, 2.6130720, 2.8213399, -1.8063687, -2.0326487, 1.1890796, -2.3557716, -2.3038208, 0.4210865, 1.4233076, -0.9454181, 2.4489761, -2.0733211, 1.4534467, 0.9295102, -0.1703898, 0.7411715, -0.5512118, -2.9706419, -1.1151812, -1.3678025, -2.3598257, 0.5751265, 2.6756483, 1.3153572, 1.6328983, -2.0480575, -1.6665178, 2.1822098, 0.0695314, -1.4384309, 0.9443320, 1.4484479, 1.0248450, -2.8508544, 0.2341084, -1.4213949, 1.6559253, -0.8073857, 0.6489826, 0.2933748, -1.6954631, 0.6207783, -2.8809275, 1.3347675, 2.8918778, -0.9212849, 1.9808599, -2.3486344, -0.7533855, 1.6153966, -0.7040993, -1.4889262, 0.1902341, -1.4720042, -2.9595362, -2.0956040, -2.5171454, 2.4648030, 2.3714531, -2.7527938, 2.7271588, 2.4627214, 0.2037258, -1.9877752, -0.4607471, 2.3585158, 2.5731924, 2.8364264, -0.4136047, -2.4475254, 2.2003918, -0.4153546, -1.7928760, -0.4486533, -1.4599542, 0.6330194, -1.7896520, 1.5765441, -2.0390398, -2.2682912, 2.8863438, -0.9739983, 2.0467034, -1.8327011, 2.0606666, -1.7197677, 0.0993556, 2.2129525, -0.3509682, 1.8160372, 0.4954852, 1.9156148, -0.7407208, 1.0864688, 0.1146062, 0.7212109, 0.4668934, -1.4117507, 1.5233695, 2.8073248, 2.0841355, -1.4175660, 2.1036003, -0.4552449, 1.5113862, -0.4480577, -0.0372429, -0.0266568, 1.3661316, 1.8626270, -0.6158325, 0.5411725, 0.7954879, -1.4862972, -2.8870824, -1.4966158, 0.8757535, -0.6525534, 1.5340295, 1.9944735, -1.0204950, -2.0404433, 1.2695190, 0.0567249, 1.6866258, 2.8222739, 1.7270615, -0.3335704, 1.7894004, -0.4064202, -2.1240006, -1.2952731, 2.2703464, -0.0481971, -0.7663352, -0.9829467, -0.3618571, 1.3486961, 0.9068771, -2.1953134, 1.6179520, -1.1793492, 0.9992519, -2.9980540, -1.8096699, 2.6668268, 2.2170685, 2.0784398, -2.4631588, -2.5356876, 0.0495929, 1.1626208, -0.5336481, -1.8412260, -1.8053093, -2.4500523, 1.7317133, 0.0107983, 2.7391192, 0.1514892, -1.2568791, -0.6559258, 0.3653213, -2.2177105, 1.3536569, 0.2658232, -1.9736597, 1.7844336, 2.5265084, -0.7032721, 2.7693546, -2.2523238, -2.3101433, -1.0563702, 2.6246571, 1.3836790, 1.0077759, 2.5375918, 2.7915652, 0.8503419, -2.4495535, 1.7738356, 0.0278383, 2.8394783, -1.9413236, 2.8525140, 2.1854173, 2.8489713, -2.4992882, 0.7992070, 2.1992675, 0.5179490, 1.0028089, 1.7632486, -1.5220355, -0.3301891, 2.7011406, 1.5002385, -2.0506836, 2.0736972, 2.3915819, 2.2062307, -0.9909251, 0.6739362, 1.9973283, -1.7055666, 1.5244390, 1.2724493, -0.7369241, 1.0076629, -0.5811846, -0.8367702, 2.4416889, 2.0333164, -2.2444115, 1.4299210, -0.6647477, 0.4234255, 2.2677747, -2.3871663, 1.2977775, 2.4722041, -1.8542578, 1.9440753, 1.3928276, -1.5132820, -0.3251049, 0.2293014, 2.9619724, 1.9695505, -1.0224292, 0.2530597, -2.2638177, 0.4565820, -2.3917006, 1.2880333, 0.3112784, -0.1088821, 1.8873471, -0.1626291, 0.1948274, 2.1001483, -2.9684215, 0.4334059, -2.3535044, -1.0716345, 1.7507712, -0.9049937, -1.6094089, -0.4239538, 2.5073730, -2.6752521, -2.1588688, -0.0555527, -0.7502794, -0.5761481, -2.9728360, 2.9298579, 2.9067315, -0.3811861, 0.5413791, -2.5651930, 2.0886722, -0.1245017, 2.6158383, 0.8308446, 0.0340583, 0.4797064, 1.7070528, -1.1513688, 0.0751017, 2.4876407, 1.6622451, -1.0804908, -1.4598348, -0.2691731, 2.9293798, 2.6897117, -0.8886027, 2.9419400, -0.9385104, 0.6015297, 1.0439833, -2.5188719, 2.4205818, 2.8157434, -2.1024495, 0.1612830, 2.3679417, -2.4781134, 2.1616249, 2.1566864, 1.8387875, 1.7152239, 0.1110830, 2.5641712, 1.5273159, -1.2843280, 2.4272793, 0.0444974, 0.8439348, -0.1591262, -2.9349659, 0.9590846, 0.2196299, 1.1397053, 1.8874741, -0.8798457, 1.5623573, -0.0895633, -2.5614916, 2.6656957, 0.0434939, -0.8197355, 1.2766194, -2.2187899, 2.2790572, -1.9150486, -0.9155493, -1.4510843, 0.1155574, 1.0969185, 2.8109355, -1.7234641, -0.1318300, -2.6500492, 2.8653438, -0.4184206, -2.2645655, 2.6972484, -1.7551477, 2.6003925, -0.5330480, 0.7380347, -2.7597856, 1.5535183, -0.4770811, -1.1093857, 0.5948248, -0.4687272, 1.8411452, 1.7587767, -1.0927595, 2.8640290, -2.3098458, 1.8663863, 1.5862325, 0.1314125, 1.0458536, -0.7646172, -1.0819508, -2.9845605, -0.6040542, -1.3812264, -0.8590106, -0.4792935, -1.6007468, 2.0735688, 1.4227639, 2.4605627, -2.5042764, -2.8835098, 1.3172864, -0.0250193, -2.8775368, -0.4255608, 2.3543043, 2.0100477, -1.5781504, -0.5336870, 2.1567110, -1.7045398, 1.9546551, 0.9515506, 0.7345600, 0.4688085, -2.2137243, 0.2085732, -1.8093718, 0.6801045, -1.7993297, -1.6959480, -2.8909550, 1.1095326, -2.7932191, 2.9436250, -2.9492451, -2.9115207, 2.8306491, -2.9910282, 0.2706203, 2.4963640, -1.5409995, 2.9202610, 0.1442234, -0.7192558, 2.9624503, 1.2237070, -1.3805099, 1.9308318, -2.5742620, -0.6461069, -1.2383225, -0.8778355, -0.8040358, 2.1966422, -1.9496062, -1.0743894, 0.9736659, 1.3239327, -2.2980897, -2.5477457, -2.6746683, -0.1941148, 1.0004030, -2.4805197, -0.9914111, 0.3951345, 0.8205907, 0.2909370, -2.3126849, -0.1780103, 1.1922563, -0.6516173, 2.6528078, 2.5947481, 1.6514745, 1.7321550, -0.9169992, -1.7754993, -2.8788090, 2.2257112, -1.7281404, -1.0265392, -1.2041813, -1.8904935, -2.6581046, 2.2612170, 1.6126237, 2.1929184, 0.9782296, 2.2771411, -2.2616154, 0.5820982, 1.5556003, -0.3174477, 1.8294926, 2.3959185, 1.4380743, -1.0364938, -0.5612529, -2.7241506, -1.3608281, 0.1252510, -1.1368598, -1.8859593, -2.6779771, 1.3544042, 2.3009793, 0.9673788, -0.6873642, 2.7019806, 0.2827624, -1.4741871, -0.1194312, 1.7083879, -2.6627625, 1.8253402, 2.7752011, 2.9310838, -1.1503875, -1.4238742, -1.6945817, -0.6421786, 2.5537171, -0.0525592, 2.3182816, -2.2303314, 1.0480174, -0.0889172, -1.7569883, 0.7820538, 1.6511023, -0.8446250, -2.3700577, 1.4099825, 0.2602278, -1.7595038, 0.3421437, 1.5854023, -1.4286550, 0.2889513, -2.2807436, 2.3066894, -0.8308948, -2.6318487, -1.5704770, 1.5268387, 1.2351520, -0.0235051, 1.0799067, -2.9780944, 0.3916404, -0.4949188, -0.9808332, 0.1837010, 1.5185750, 1.5823746, 1.5232917, 0.0610893, -2.3421017, 1.3094164, -2.8547603, 0.2053670, -1.7366316, -1.6636797, -1.6752903, -0.7232966, -0.9318375, 2.9528376, -0.8717759, -1.5211502, -0.3874390, -1.7523671, -1.7500350, -2.6141488, 2.0759522, 0.5868125, -2.9356857, 1.5128899, -0.6578224, 0.1554613, -1.8638711, -2.5030703, -1.6118951, 1.8279723, -0.3803986, 1.0331197, -1.3796464, 1.3119082, 2.5381730, 1.7136926, 0.4799174, 1.4264906, 0.6885764, -1.9415673, 2.5760695, 1.7399748, -1.6398179, -1.7068777, -1.9607567, -0.8467240, -1.0308238, 2.2977166, 0.7525824, -1.2507189, 2.9568788, 1.2112083, 0.7690835, -0.7898136, 1.8817608, 1.7913914, 0.2251665, -0.6059082, -1.9139421, 2.2127751, 1.4361557, 0.8357342, -2.8524577, 1.4986006, -0.5953462, -2.9363473, 0.0606835, -0.0385475, -0.0208070, -0.5249525, -0.2976299, -2.8288430, -0.7195562, 2.9201880, 1.3438886, -2.5027139, 0.2439483, 1.3399691, -2.7525528, 0.3276044, 1.5041122, -2.6484086, -1.5322018, -2.5770106, 1.8416803, 2.9047453, -1.0825098, -0.6452352, 2.6939686, 2.9244394, -2.6393954, 2.4005253, 1.4099729, -1.0819270, 2.2677605, 1.8017315, -2.6714056, 1.2796746, -0.8757883, 2.5600538, -1.5163289, 0.6771283, 1.8185592, 2.9784332, 0.9053742, -0.4313803, -1.8000428, -1.3621711, 2.1645309, 0.8445679, 1.2326859, -2.6560554, 2.7602635, -1.1627106, -0.8962695, -2.7193658, -2.6728740, -1.0947077, 2.5415077, -0.6208173, 1.9773604, 2.6974809, 2.3587526, 1.7432664, -1.2625170, 1.5554567, 1.4845742, 2.2335124, 1.3361048, -2.2743757, 2.3466601, -2.9508771, -2.5506686, -1.6735927, -0.1226048, -2.4126001, -2.8554716, 0.6305935, -1.9387754, 2.2218518, -0.3987674, 2.6159853, -2.6609471, -0.1377921, -1.5580009, -2.3826540, -2.3703519, -1.0360915, -0.8030908, -2.4410728, -0.4246388, 1.2314991, -2.1234546, -2.0944902, -2.9210669, 0.2224948, 1.4488822, -1.9298921, -0.2932189, -1.2345913, -0.7871992, 1.0550294, -0.9689441, 2.5735760, -2.2457420, -0.2531746, -2.7646142, -2.6662199, -1.4601966, 0.1533270, 1.7021413, 0.9304762, 0.5342932, 2.4561644, -1.9401211, 0.6946785, -1.4425679, -2.5583503, -0.6560180, -0.0241282, 1.8503818, 2.2189686, -0.3699883, -1.8403735, 2.6309801, 2.6467524, 0.2294531, -2.2783243, -0.8389042, 0.9790286, 2.5188409, -1.7929783, 2.3838328, 0.5797630, 0.0871403, -0.4365213, -2.3517911, -2.2851528, 2.4828311, -2.8675854, 2.0439084, 2.2227963, -2.4083532, 1.5754750, -0.7711952, -0.0089817, -1.5843608, 1.7598023, 1.9227750, 1.9241869, -1.7320216, -1.5012929, -2.1788065, 2.1266690, 2.3677150, -2.6678122, 2.3896712, 2.8317094, 2.8103928, 0.1462804, 1.3920639, 2.5270530, 0.4068558, 2.7432884, -2.8560098, -0.7954787, -0.6188917, -1.5747237, -1.3472437, 1.1992764, 1.7229445, -0.7777533, 0.5697030, -2.2059627, -0.1206169, 2.7484155, 2.5150860, 1.4161554, -0.3554038, 0.5712984, -2.0228476, 1.1048671, -2.3724504, -1.9932279, 1.4108035, -0.8369163, 0.7281219, 1.9145712, -0.7517635, 2.5360429, 0.3952076, 0.1384339, -1.5711084, -1.0475017, -2.8993824, 0.2294581, 1.7702190, -1.7855732, -1.7244854, 2.9805645, 1.8084436, 1.4618432, 2.1803009, 0.0368244, -1.7283191, 2.3465789, -1.8633881, 1.9126210, 2.7649008, -0.7919891, -0.4859682, -0.8054771, -1.6987411, -1.4609200, 0.6053015, -0.7506624, 1.2947618, 1.1232559, 1.1270402, 2.6973879, 1.8038153, -0.5751921, -1.2583240, 0.0904762, 0.4308282, 0.4732877, 0.9925409, -0.0152690, 2.6041520, -1.1899474, -1.3147278, 1.0895998, -2.5747954, -0.9394877, -1.8694715, 0.8817487, 2.3171523, -2.0790480, 0.3750969, -2.2346834, -2.2474153, -0.2756334, -2.7842666, -0.0816610, -0.1475642, 2.7035054, 0.8336616, 0.4984691, -0.4854758, -0.2341211, 2.0129353, -0.0660161, 2.2114884, 0.3037827, 1.9673423, -2.2380088, 1.4223075, 1.8099028, -0.0678707, 1.5786408, 0.0108818, -1.1576123, 1.1265618, -1.9881813, 0.8473715, 2.0129072, 0.2173467, 2.0542079, 0.0164830, 2.7729896, 2.3325292, -2.2043484, 1.8379370, 2.1201610, 1.2277867, -0.7788619, 1.9693307, 1.3584365, -0.1497266, -2.1225370, 0.1134772, 2.4487096, -1.2179779, 0.1022956, 0.4022882, 0.6778478, -2.0045123, -2.7266015, -1.5250371, -2.3761375, -1.1647113, -1.9563275, -0.1562890, 0.2076763, -1.1455079, -2.8717092, 0.4819850, -2.9070120, 1.6693169, -0.2535900, -1.5920682, 1.2585261, -2.7653194, -0.7283021, 1.6258913, 0.5944252, 0.9091932, -2.4473209, 1.3018897, 2.0950228, 1.6571828, -0.4970854, 0.1944918, -0.2046651, 1.1827076, 1.2771377, 2.4153309, -1.9008987, 1.5186582, -2.8042124, -0.5931141, 2.8437587, 2.1218702, -0.4198787, 2.1713236, -1.8087616, -2.2683743, -0.9411735, 2.6870569, 1.4497146, -1.1804663, 1.9932495, 0.3149791, 1.0719744, 0.0984482, -2.6647460, 2.2269163, 1.5884002, -0.6567368, -1.0235776, -1.8693938, -2.6308216, 2.6819636, -1.3878753, 0.9302169, -1.5337079, -0.5788498, -1.1555926, -1.0434161, 1.7731074, 0.3433668, 0.3063468, -1.6635083, -1.7532285, -0.7955938, 2.3394021, 2.7878534, -2.2605512, -1.7922730, 2.7203636, -0.9621021, -2.1921803, 1.2195527, 2.8806688, -2.4915450, 2.8369375, 2.5636676, -1.4214774, -1.7461559, -0.7285992, 1.6627471, 2.1181658, 0.4761422, -1.5442654, -1.6698167, 2.9793307, -1.7171737, -2.4075884, 2.0151543, -1.4545768, -1.1230040, 2.0499649, -1.4095920, 2.0825583, 2.3892901, -2.0336644, -0.0118636, 1.8749410, 2.0440656, -0.5109799, -2.7895908, 0.8674895, 1.6403507, 1.8592649, -2.1421364, 2.2766556, -2.1186914, -0.1599779, -1.2398866, -1.0256814, -0.6780169, -1.9341863, 2.8667835, -1.1645547, 1.3479208, 2.3497351, -1.8430091, -2.4289114, 0.3794579, 2.1760173, 2.1181415, -2.0198784, 0.3510489, 0.6952729, -2.5110484, -2.6876718, 0.0395676, -2.6922106, -2.5189703, -0.2205209, -0.2177776, 2.1239582, -2.7422506, 1.8533318, -1.5491771, -2.2096469, -0.7562984, -2.2637651, 1.6841832, 1.7383742, -1.6589949, -2.5038076, -0.2615316, -1.9309739, 0.8423034, -1.4666704, -2.1967402, 2.1292362, -1.9081907, -1.9814837, -0.8253889, -2.9021205, 0.8199907, -2.0003912, 0.1376921, -0.5368703, 0.0750305, -0.3065416, 0.3092508, -0.0178791, 1.4467565, 1.0653375, -0.6588741, 2.2663508, -1.3065324, -1.6360253, 2.8210452, 1.7020409, -1.5406240, -0.1684521, -1.0389903, -2.9130172, -1.4474368, 1.3379879, 1.6903393, -2.8828161, 1.2478730, -0.4587459, -0.9469120, 1.3073762, 0.5852810, -0.5553216, 2.6110151, 2.5375500, 2.9969520, 2.5805498, 2.5097631, -2.4489935, 0.3736490, -1.8861671, 0.4797075, -0.1096499, 0.5951288, -2.2638333, 0.2162072, -0.4662941, 1.0594802, 1.0441492, 0.6554590, -2.4261722, -1.7994654, 0.8768931, -2.4375670, 0.9620192, 2.1888203, 0.2353364, 1.7287926, 2.6356950, -0.9026702, -2.5609485, 0.5887544, -0.0239319, -2.7719913, 2.7195631, 2.0416362, 2.5459319, 1.6045233, 2.9663797, -2.8016864, -2.3523623, -0.4215878, -1.0718383, 2.0998721, 1.5301210, 2.1176727, -2.7780391, 1.7286120, -2.6241603, 0.3906998, 0.4807556, 1.0679425, 2.3459295, 0.1510823, -1.7085780, 0.0904466, -1.9337564, 1.5140194, -1.7628954, -2.3811007, 2.2018491, 2.8487460, -2.0050358, -2.2005021, 2.5112441, -0.7223938, 1.0701171, 2.5105630, -2.7951292, 2.2313628, -2.1720439, -2.1883086, 0.2667828, 1.8538338, -2.4452625, 0.2954414, -1.3296695, -0.2395499, 0.3546013, 0.0421279, 2.2640704, -0.9156372, -0.5531985, -2.1071361, 2.9982349, -2.1981827, 2.5677621, 0.4827933, -1.4028493, -1.0334567, -1.1902379, 2.6360568, 2.3873285, 1.0488301, 0.1375960, -0.9205618, -0.9563852, 1.9676478, 2.7275016, 1.3211527, 2.4861491, 2.1786119, 2.2025499, 1.8303168, 2.6688862, -1.6750502, -0.2464646, -1.0835387, -2.8926639, 2.6566081, 2.6577941, 1.2603045, -2.7018988, -2.1712392, -0.9674072, 1.5192056, 2.7520007, 1.2181005, -1.6150628, 0.8751712, 1.2648879, 2.0925492, -0.4581662, 2.4874782, -1.7133415, -2.2969536, -2.7243853, -1.7411121, -1.0301318, 0.4247473, 1.5254091, -1.9301725, -2.4502599, 0.2472917, -1.9197811, -2.2296162, -1.7509368, -1.7915150, -0.5346179, -1.3637693, -2.4848755, -0.5684317, -0.6001913, 2.0430571, 2.1770603, -0.3459084, -1.8985652, 0.1640965, 1.2134146, 0.3903754, -2.8831126, -1.3273170, -0.2779266, -0.6204053, -2.5187881, -0.3064017, -2.5926724, -2.1757831, 0.7774078, -0.4810295, -0.8857999, -2.1970970, -0.6876810, 1.2120541, 0.8681101, 1.0048784, -2.9791566, 2.3956318, -1.4502999, 1.3146367, 1.0799829, -0.0530063, 0.7909867, -1.5148820, -0.9434765, 2.2066131, 2.8334078, 2.1163058, 0.7583675, -2.2338394, 1.2552310, 1.9976220, 2.0550137, -0.3278553, 2.3764718, 0.0716276, -2.6261811, 2.7710924, 1.0232403, 2.1647121, 2.3160377, 0.8786910, 0.9762209, 2.0562598, 2.8689821, 1.7097367, -0.2276635, -2.0843820, 1.5413729, 1.2144184, 2.3445054, -1.3333976, 2.3542553, 1.9507573, -2.0846381, -0.8822907, -1.5897957, -2.3743079, 1.6269784, -0.1624662, 1.4089913, -0.6866656, -0.1026869, -0.4627415, 0.4376914, -2.2811183, 2.7746025, 1.9024182, 1.8305045, -2.3894669, -1.1320691, 0.1273308, -1.8920031, -2.1072826, 2.8710650, 0.5926710, -1.6945915, 0.6744432, 1.6546728, -2.7324297, -0.2784905, -0.0396806, 2.2989942, 0.4492955, 2.5024597, -2.3844897, 1.3639201, 0.7796929, 2.1911249, 1.6153481, 2.5959739, -2.2786338, -0.9713121, -0.6678350, -2.7097033, -1.2516116, 2.0754631, -2.9541450, 0.7010578, 1.0594508, -0.8029203, -2.5864872, -2.4297462, 1.9708300, 2.0835319, -0.1583538, -1.8530892, 1.3380589, 2.1516623, 2.9037409, 0.0622603, 0.3881647, -0.7544381, -0.8699020, 1.2830923, 0.1492592, -1.5860480, 0.6063964, 2.4147003, -1.3590892, 2.4634768, 2.4261216, -2.4873523, -2.1918746, -1.5925929, 0.9976562, 1.3488293, -2.2870478, -0.7446022, -0.5045668, 2.7000690, -1.5730242, 0.5090217, -1.5719353, 1.3733943, -1.3629190, -2.7166084, -2.6699432, -2.5257622, 1.2646208, 2.0264385, 2.1829318, -1.9033099, -2.6862746, -0.2514949, -2.8146252, 0.8767729, 0.5471455, -2.6696753, 0.0272890, 2.4731126, 0.7999632, -0.9398487, 2.4353800, 2.8749091, -1.5352026, 1.7176044, 0.0257038, 1.9524180, -1.6936977, 1.7043370, 1.3907389, 0.2048890, -1.5076441, -1.9342734, -2.7820873, 0.6639610, -2.3845930, 2.9769954, -2.5113591, -0.5793763, 0.0886797, 0.9808831, -0.3785050, 0.3401570, 1.7641522, 2.6898115, -1.2470103, 1.2761258, -0.3294719, 1.7726404, -0.7499842, 1.6921753, 0.6398271, 2.4651193, 0.1981076, 1.9038489, -2.7441410, -0.1513170, -1.1758892, 2.3489635, -0.1305970, -1.2767934, -1.4923082, 0.2499852, -2.3128284, 2.9616162, 0.4069864, 1.2262765, -1.3376729, -2.3466358, 0.2113706, -1.2525789, 2.1794118, 0.7609708, 1.1058286, -2.6200083, 1.2087975, -0.5480926, -1.9493777, -0.1925285, 0.8909709, -2.9261262, -2.1813570, 0.5978792, -1.9435208, -0.6738217, 1.3456709, -1.9538264, 2.1235054, 0.7846748, -0.9568173, -0.4575311, 0.9139543, 2.6015249, 0.9105580, 1.5828172, -2.5057796, 0.1690734, -2.7834854, -1.1476718, -1.8705579, -2.8723490, 0.1594225, 0.2372246, 1.4897073, 2.1790878, 0.3062226, -1.4595287, 0.5553393, 2.7690421, 2.4160789, -2.1611479, 2.0662809, -0.0503450, 1.5794443, 0.1496704, -0.0461467, 0.5927543, 1.1243584, 2.7320693, 1.8223024, -1.8444968, 2.0461778, 1.6754487, -1.3348045, -0.1815448, -1.5853427, -2.2731073, -2.1044791, 0.1053112, 0.1613209, 0.5947929, -0.3741569, 0.3398675, -1.2797373, 2.8370799, -2.7579305, -0.5371945, 2.4338530, -1.7262093, 2.9887283, 0.6611854, -2.6503980, 2.8344812, -1.1951997, -2.5178830, -2.9407812, -1.5775381, -1.3306149, -0.3496602, -2.9885064, -2.9742128, 0.2768614, -0.6552048, -2.5785971, -1.8363719, 1.9432255, 1.0619350, 0.5770033, -2.7492435, -1.1177075, 1.8683854, 2.6601875, 0.5911520, -1.9301417, -2.2200610, -2.3763833, 0.7509133, 2.8127188, -2.7672291, -1.9257706, -1.7144899, 0.3417885, -1.0503140, 0.3706718, 2.7087407, 2.8257293, -0.2023477, 1.1021840, 2.6273272, -2.1947236, -0.3813788, -1.4020156, -2.1764302, 0.6045280, 2.3070371, 1.6144006, -1.1072205, -2.1302665, -1.3946419, 1.6292418, -2.0361439, -1.3361644, 0.4697154, 2.5837744, 1.8095259, 1.1774035, -0.6499685, -2.8780525, 1.1507646, -1.4859503, 0.3552076, 2.8276401, -2.0880110, -1.7843252, -2.0325906, -2.3015894, -1.0655150, -2.3076659, -0.3614350, 1.1051697, 1.7574827, -0.1120807, -2.7035493, 0.8245853, -2.3934296, 2.6660415, 1.1473352, -2.9703491, -0.8007502, -0.0644438, -0.1961591, -1.8772072, 1.5433241, -0.5385926, -1.4212797, -1.0211238, -0.1551940, 0.8031688, -2.9288906, -2.6721367, -1.8534217, -0.3704660, -2.0248473, 0.2870531, 2.0068995, -0.3743794, 1.5379989, 1.6324375, 1.0971755, 1.5737097, -0.3293832, -1.3214089, 1.8083159, 1.7741964, -1.2373244, 2.3411707, -1.8500467, 2.2338612, 0.3290070, 2.0325508, -2.4686503, -0.9197652, -0.2144817, -2.2833099, 0.5692197, 2.6960850, 2.1683006, -2.5987084, 2.2681497, -2.6014233, -1.9968006, -0.4116551, 2.6450597, -1.8897782, -2.1456941, 0.5601458, -1.4572547, 2.4945931, -0.5890768, 1.0158279, -2.7261335, -0.4221739, -0.3096224, 0.6284411, -0.1357548, 1.7322773, -2.5577764, -2.0866254, 1.8967980, 1.1772880, -1.2552277, 1.7320554, -0.5635451, -1.7635551, 0.4161167, -2.8751811, -2.0859857, -2.8448780, -0.5638894, -2.5845313, 1.3298291, -0.0995864, -0.7437871, -1.5134011, 0.4697774, -2.0840665, 1.0768697, 1.1095175, 2.3561757, 1.3246956, 1.4298004, -1.5169908, 0.0360828, -2.2263907, -1.2710197, 0.2151140, 2.4815174, 1.4056828, 2.6365637, -0.4000702, 2.6677752, -2.1006880, 2.8545175, 2.6294130, 2.2666902, -2.2537960, -1.3387168, -2.8420489, 1.1106914, -0.3617431, -1.6405591, -1.8032141, -0.5758951, -1.4171396, -2.4826411, 1.9993781, -2.9416468, -1.6624572, -0.2203050, 1.8744349, 1.1213904, -2.2237631, -0.3181067, -1.7737564, 2.1686627, -1.9774541, 1.5600586, 2.2319455, -0.0206276, 1.0902685, 0.1406664, -2.3964215, -1.0701506, 2.5274463, -2.6133460, -2.1614065, -1.1247959, -2.4911528, 2.9510151, 1.7087676, -1.5884239, 2.0606670, -0.8213677, -2.5799532, -1.3870779, -2.4475699, -1.3209841, -2.7539764, -2.3049394, -1.3143030, 2.0756815, -0.3019429, -2.4794452, 0.9942203, -1.8081423, -2.9752720, 2.6501789, -1.5832222, 1.0636093, -1.7494094, 0.0426915, -0.4736353, 0.7804029, 0.9621360, -2.4497495, 0.2741319, 1.9975180, -1.3295768, 2.0010891, -1.7120305, -2.5347273, -2.8669229, 2.3787626, -0.7728482, -2.3643162, 0.6151539, -0.5374066, -0.7053683, -1.2250020, -2.1119322, 1.3864097, 2.1404985, -2.2664866, 1.3658068, 2.4336304, -1.1875248, -0.7889532, 0.4601722, -1.4412435, 0.0906771, -1.9964797, -2.5196145, -0.1917852, -0.8596172, 2.1936717, -2.5423501, -2.3216182, -1.2585074, 1.3162487, 2.3324735, 2.1856908, -0.8834977, -2.8425735, -1.0127533, 1.9236920, -2.7994454, -1.3270982, 0.7768564, -1.9756597, 1.6298986, -2.4832723, 1.7647925, -1.6345474, 1.0022133, -1.1905982, 0.7457897, 2.7429837, 1.9759582, -1.6607056, -1.9702077, -1.6373902, 2.6224172, 0.9900805, -1.2477478, -2.6220020, -1.1326395, -1.3428861, -2.3558839, -2.7903751, 2.5246591, 0.7783886, 2.8879846, 0.9432319, -1.5228673, 2.4896710, -1.6913283, -2.0518800, 1.2474727, 2.6826994, -1.2731229, 2.6963761, 2.3802032, 1.7117208, 2.9542152, 2.3170798, 0.4658717, -2.2405910, -2.8058879, 1.3326676, 1.5604391, 2.9890944, -0.9824073, -1.1957598, 2.9174865, 2.7830808, -2.0121675, -0.3425043, 2.1806841, -2.5282988, 1.4721568, 1.5858297, 2.3531799, -1.6966190, 0.6160430, 1.3133434, 1.5853973, -1.5977095, 0.8816517, -0.9978255, 2.3068120, -1.7157946, -1.6666831, -1.4251991, 2.6907201, -0.4827803, -1.4346963, -0.6282592, 0.1205402, 2.3141665, 2.7658952, -0.6884616, -1.9647709, -0.8059191, 2.9633826, -1.1983466, -2.8369729, -0.9915246, -2.9122215, -1.4598525, 1.4251226, -1.2202495, 1.7604875, 1.0537018, 0.2518215, 0.2831879, 0.4888529, -0.0793024, -2.1938895, 0.1239677, -1.3362001, -1.8578248, 0.4351783, -2.9960388, 2.1991783, 1.9312510, 0.2113810, -1.7473689, -1.7230323, -2.8925409, -0.2849319, -1.7365814, 1.4448850, 0.6010296, 0.0821969, -1.8729027, -0.9417042, 0.1364363, -0.9591691, 0.3936291, 1.9329972, -1.9931972, -2.5920792, 2.6290024, -0.9432626, -1.5159444, 0.4074028, 2.5730582, 1.8909976, -0.1442841, 1.9008030, -1.3268289, -1.1818113, -1.4560150, 2.2867319, -2.6360575, -0.4078153, 0.6478640, -0.4965201, 0.2024884, 2.4958319, 0.0878892, -1.1460084, -2.9895517, -0.4838701, -1.6463294, 1.3392489, -0.2977795, 1.0958657, 0.5749929, -2.7072317, 2.6020219, -0.8543875, -1.8765973, -1.6382005, 1.8668931, -1.0873452, -2.7504543, -1.4513439, -1.6393104, 1.0409971, -1.2371563, -0.8731796, -0.2202245, -2.2300223, -2.9356570, 0.1469985, 0.2818056, -2.8745030, -2.1715993, 1.1699482, 1.8355247, 1.3912570, 0.5058712, -0.8916854, -0.4915113, 1.0460356, 1.2335263, 0.7296297, 2.1511645, 2.8714593, -1.5910806, 0.5589097, -0.9858860, -0.6015005, 1.9779208, 1.8344687, 0.1007509, -2.2146005, -1.3824019, -1.2401719, 2.5509225, 1.8380428, 0.8735180, -2.6764537, 2.0708595, 2.2006384, -1.9936738, 2.3215863, 0.5550796, 1.3622842, 1.5582998, -2.6944466, 2.0657482, 1.2281495, -2.0411221, 0.1551947, -2.1569098, -1.9515764, -2.8931522, -0.6143356, -2.8586871, 2.1344645, 1.5027904, -1.1320093, -1.9069605, -2.3865469, 0.0865800, -2.2625362, 2.5061309, -2.1300191, -0.8228554, 1.7100123, -2.5504072, 1.4737917, 0.6860185, 1.7332712, 1.1635342, -1.0954927, 0.3642095, -2.4796275, -2.5708831, 1.7098098, 1.2750384, -2.4489841, 0.9968452, -0.2344247, 2.1598739, -2.1296320, 1.2849730, 2.9004492, -0.4249450, 2.9694132, -0.6214346, -2.1356312, 1.6012182, -2.4802022, -0.7490786, 0.2968970, -0.2617875, -2.4374431, 0.1976074, -0.4421949, 0.9881528, -0.0979232, 0.9194813, 2.1372353, -0.9596431, 2.9142996, -0.5905128, -1.6692299, 0.1172650, 2.4803394, -1.1399013, 1.0105139, 2.3048271, -0.5220126, -1.5756474, 0.3989916, 1.4583711, -2.0252435, 1.1893807, 2.8674617, 0.6006032, -0.2544153, -1.7553188, -1.5826904, 1.5985447, -0.9667816, -2.9356215, -2.0779634, -2.1053824, 2.0617861, -2.7177271, -1.9723303, 2.2749727, -0.2408216, -0.3456665, -0.4287933, -1.6367401, 1.3440039, -1.4285780, 0.9988543, 2.5675404, -0.9350083, 0.3689639, -0.7772942, -2.6024307, 0.1977350, -2.0341483, -0.9231166, -2.8147969, -2.3710620, 1.4148699, -1.0040100, 1.6424507, -1.4341628, -0.8580631, -2.4266245, -2.1105005, 2.4898354, 2.3359867, -2.5630399, -2.6789204, 1.9127934, -0.1141182, -0.5588759, -0.4348335, -2.9541023, -2.5195122, 0.2682207, 2.2342001, -0.0144419, -0.2828619, 0.5806094, -1.8649623, 0.1044442, 0.1718160, 0.5690955, -0.8789714, -2.1380722, -2.0781667, 1.1598245, -0.7122917, 1.3703097, -1.6395478, 1.6750340, 0.8670001, -0.7514901, 2.0820957, 0.5630420, -0.3255491, 0.1307405, 0.3578978, 1.2537464, -1.6350996, 0.6377541, -0.5358448, 0.4217854, -1.6290824, 0.8403094, -0.2316662, 1.7062377, -2.5142928, 2.0408486, -0.1151093, -0.0437346, 1.0053876, -1.8123590, -1.5629364, 1.0033834, 2.9603801, 1.9759039, -2.1909321, -1.8000945, -1.8033442, 1.7886091, 2.8590835, 1.7507013, 1.8628638, -0.4048354, 2.3498062, 1.2534404, 0.7666865, 0.7767260, -2.7815885, 0.1246048, -2.1483778, -1.4876883, 1.4951553, 1.7687766, 2.1899270, -2.8363435, -2.1401767, -0.2196199, -1.6967072, 0.0640728, 2.8603658, -2.2061854, 1.8528339, 0.7894653, -0.7506829, -2.4693573, 2.1301080, 1.0546223, -0.0962793, -1.9755802, 0.9323166, -1.9334487, 1.6642278, -0.9410379, -1.3393376, 2.0902843, -1.1949574, -2.3690436, 2.0585375, 2.3431140, 2.1646507, -2.0852736, 2.9147199, -2.2847582, 0.8399278, -0.4146832, 1.8667618, -1.2460347, -2.4020539, -1.7901324, 1.4619975, 0.5443307, 0.8602715, 1.4287787, -2.4070451, 2.9041473, -1.7367635, 0.2297257, 1.4885590, -1.2640421, 2.6972748, 1.5321458, 1.9553417, 2.0705884, 2.4547643, -1.3894104, -2.4259533, -0.6708968, -1.9540437, 0.6347054, 1.3335254, -0.0653491, -2.5887835, 2.4348541, 1.5460638, 1.2032513, -1.8023726, -1.8156116, 2.7115496, -2.3824459, -0.9364422, 1.4892841, 1.8382299, -0.5969594, 0.7445086, 1.4548807, 1.4986223, -1.8914061, 0.9543085, 2.3452856, 2.0844116, 0.3362636, 0.3266029, 2.5326227, -2.7692902, 2.1274446, 1.4189904, 2.0113447, -2.2924027, 1.9789362, -0.8489214, 0.0032110, 0.5386044, 1.4569338, 0.4161098, -1.3646930, -0.5256376, -0.9341384, -0.7707897, 0.7397591, 2.9634760, 0.7835688, 1.4457069, -2.3991822, 1.1802661, 0.3599966, -0.3807637, -0.9741455, 0.8160572, 0.7545990, 1.5281221, -1.7064102, 2.3145798, 0.4138967, 0.0080878, 1.7316596, -0.1906212, 0.9856518, 1.8017505, 1.0753052, 2.6884464, 1.3334587, 1.7163678, 2.1753337, 1.0540864, 0.2632724, 2.1843094, -0.0189843, 1.6749856, -2.0769146, -2.0023542, 2.2079456, 1.4343978, -0.4863993, -2.3545898, 2.2855906, 2.1382028, -0.3198186, -0.4499920, 1.4475024, 2.2209056, 0.1828206, 2.9313151, -0.5939346, 1.8858224, -0.7990744, 2.4710912, -2.5478098, 1.8537716, 2.6167086, -2.1447761, -0.5894952, 2.7082154, 1.5862656, -0.4990052, -2.0286521, 1.8722417, 0.9393662, -2.8801321, 2.6700585, 2.3419774, -1.1845118, -0.3896525, -1.6215322, 0.8564225, -0.9119907, -1.1086000, 0.9188915, -2.9143821, 1.3306744, 1.0228832, -1.9844318, 2.1462350, -2.1087871, 1.4719578, -2.5239158, 1.2374466, 2.8419042, -0.3983346, -0.9544493, 2.7741302, -2.8661975, -1.0741885, 0.9163568, -1.8355004, 2.1962671, 2.5341883, 1.9174696, 2.4535603, 1.4404258, 0.8024513, 2.8186899, -0.5122680, 1.3776595, -0.1999817, -2.4694387, -1.8423772, -0.8833461, -0.2978423, -0.6055854, -1.9466419, -0.2747254, -2.8026794, -1.3913979, 0.3874949, 0.5638977, 2.7431743, -0.3696934, 2.4944203, -0.3831454, -2.5151688, -2.7415598, -1.6991686, 1.0248417, -1.8496030, 1.3068745, -2.8831996, -0.5700131, -2.8609493, 2.4679580, -2.3265725, 2.9956260, 2.7468966, 2.1879517, -1.2588164, 1.0310607, 1.7516573, 2.3355871, 1.6707218, 0.6599345, -0.9708529, 1.0011215, -0.2882469, -2.0996034, 0.8265409, 2.2907166, 1.7994236, 2.9149945, -1.2469864, -0.4603723, -2.1175373, -0.5255891, 0.1655068, -1.8140278, 1.9789757, 2.3861471, -1.2708822, 2.9399897, 1.3741011, -0.0533968, 0.1744490, -2.2308974, 1.1352610, -1.1537208, 0.1955410, -0.0566351, -1.1705676, 2.6043634, 0.7112401, 2.8124548, -0.4428203, 0.8160651, -0.7061883, -1.8251266, 1.9906715, -2.9342624, -2.5276212, 2.8104385, -2.3560173, 0.9096217, 0.0385778, -2.3423472, -0.3470709, 1.1638747, 0.9246304, 0.2586792, -1.4162416, 2.1994784, 2.6554653, -0.6096244, -2.3305967, -2.8954436, 0.1330814, -2.7623110, 2.1394275, 1.4260773, 2.0999818, -0.1562584, 1.0664624, 0.9547899, 0.1630216, 0.9634150, 0.5034119, -2.9874824, -1.1495640, 2.6097814, 1.7888631, 1.6711598, -2.6360701, 1.3185020, 2.4130806, 2.8499430, -1.0849688, -2.0409181, -2.0036123, 2.4031092, 2.6985808, 0.6312884, -1.0233723, 2.0491135, 2.5168992, 2.1805834, 2.1919486, 1.0300175, 1.4413403, 1.2316262, 1.6077271, 1.8936122, 2.7154366, -2.6950499, -0.2600532, -1.4892618, -1.4874353, 2.0143844, -2.6478103, 2.0493756, -2.0234339, -1.5749134, -0.6159152, 2.9018064, -0.4724526, -0.1607710, 1.0310402, -2.7773242, -1.5743120, -1.6720481, -0.6231065, -0.6072798, -1.2795436, 1.6342514, 1.5008239, 2.4020245, -2.6271940, 2.8797821, 2.7083003, 0.0678311, 1.4427988, -2.4427147, -2.6708443, 2.4423590, -2.6467078, 1.0721407, -1.5707750, -2.0112446, 1.5786438, 2.5559411, 2.6470925, -0.9499886, 1.1198973, -0.9830970, -2.0395555, -1.7276013, -1.7949309, 1.7108216, -2.4965365, 1.6460105, -2.6798496, -0.7410559, 2.5064648, -2.8055096, 2.1528218, -1.4353253, -0.9761702, 1.1152755, -0.8178279, 0.4797950, -2.5587394, 0.6984237, -0.9623368, -2.6465782, 1.7435817, -1.7805823, -2.6711588, -0.6983257, -0.7785508, -0.4153079, -1.8700001, -0.5100887, 0.4892980, 0.5940482, -2.9246779, 2.7944251, -0.8256056, -1.2162793, -2.7514134, -2.0700084, 2.6734929, -2.7718990, -1.5945223, -1.6719115, -1.9673106, 0.4970367, -2.2521213, -0.6385819, -0.5873048, -1.1378776, 1.0352296, 1.4659245, -1.1016698, -0.5214768, 0.9515308, -2.2140360, 2.3508649, -0.7992391, -1.9054216, -0.6580474, 0.1606884, -0.0524904, 2.4062186, 0.1945970, -0.7424176, -0.2166471, -2.6823868, -2.5607198, 2.8247231, 2.7692395, -1.7443445, 0.3703159, -1.1699113, -2.9387700, -2.9156629, -2.5570383, 2.2215993, 2.6691318, -2.3178151, 2.5935947, 0.4973319, -1.9708060, -1.2855315, -0.4560627, 0.1388137, -0.1190655, -0.9399163, -1.0808297, -1.5195645, 1.0659751, -1.2225774, -0.0175797, 0.5847465, -1.2617767, 2.5930009, 0.8744449, 0.8295115, -0.4094404, -0.9417693, -1.5570571, 1.0777823, -0.6826838, -1.4179356, 1.7262894, -1.2775537, 2.7183604, 1.1270466, -2.4492789, -2.4486320, -2.8079784, 2.6450310, -2.3187295, -1.6442143, 0.5164891, -1.7218945, 0.8420268, 1.4848238, 0.4874570, -2.1287931, 0.0073778, -2.2592502, -1.4946602, -1.9715836, -2.9927580, -0.9756847, -0.5149461, -0.0019090, -2.4376672, -1.6995303, -2.3134671, 0.2801216, -0.8816778, 1.7102261, 1.9113002, -2.4436689, 0.1821059, 2.6820474, -0.6337975, -0.8742863, 0.4504672, -1.5976924, 1.0861471, 2.6455887, -0.1644054, -1.0618345, 2.6485422, -1.4133354, -0.0226031, 0.5506681, -2.2755938, 1.7691007, 2.4963595, -0.1895660, 1.2543061, 2.9469180, 2.0480970, 2.9886588, 1.4222513, 2.5540072, 2.5631159, -2.5521365, 1.6902883, -2.4523802, -0.6922781, 2.8193538, 1.3396464, -0.9070046, 0.7374750, -1.3973326, -0.8695349, 0.1899748, -0.5670679, 2.4539491, -0.5808583, -0.1899169, 0.5374748, 0.2474853, -0.1808849, -2.5566105, 0.5858190, 0.5751347, 1.7000901, 1.3494482, -0.3273663, -1.7690815, -0.4544222, 1.0417141, 0.4704274, -0.7775279, 1.6559064, -1.4779283, -0.3590098, -1.5145653, 0.6660043, -1.6080120, -2.1400555, -2.4795150, 0.2843529, 0.0192157, 2.1315111, -0.0062308, -1.9737522, 0.0250530, -2.4627370, 2.8519110, 1.3958408, -0.2458899, -1.7756610, 2.4407122, -0.0548962, -0.7779546, 1.3940032, 1.6705456, 0.3650630, 2.5473723, -0.7633423, -0.8294498, 2.2070422, 2.9318826, 2.9185170, -0.4793817, 1.6910870, -0.3342982, 2.4309055, -0.7859731, 1.1431083, 2.7917222, -2.1872324, 0.7902615, 2.7145713, 2.8181722, 0.3089837, -0.7565712, -0.5278929, 0.3983347, -1.7681877, -0.6720348, -1.6406751, -1.1258096, -0.4596248, -1.5472381, -1.7177256, -1.7359934, -1.2998348, 1.2397141, 2.4377745, 1.5589825, -0.1293547, 0.1145945, 2.1465410, 0.2499005, -1.9434647, -2.2660840, 1.3411908, -1.7010840, 0.3599597, -2.8917037, 2.4428361, -1.5274042, 1.5864144, 1.9509467, -1.6588264, -2.8732118, 0.2632841, -1.4830543, 1.3760142, -1.4296066, -0.3809071, -0.9663035, -2.3660569, -2.9592627, 1.2537641, 1.8778464, 2.1051714, -0.4880784, -1.9583354, -1.5032071, -1.6671394, 0.3507568, -1.5467153, -1.3937717, 1.9309353, 0.6404032, 1.5306217, 1.5217275, -2.4304550, 2.1690436, 0.2565965, -0.0422210, 2.9900164, -1.9088071, 1.8526882, -0.5216945, 1.8002666, 2.5324674, 0.7385079, 0.0404383, 1.1827051, 1.6380245, 0.5772310, -0.1868728, 2.1702435, 2.5003389, 1.3660395, -2.0420723, 2.7540333, 0.7169311, 0.2392530, -2.0502345, 0.8596064, -1.4551128, 2.2499805, 2.4229660, -1.9509252, -0.9747925, -0.4837853, -1.2428590, 0.3776809, 2.1170021, -0.6560022, 0.0190591, 2.2737589, -2.6147676, 1.4997610, -2.8825514, -2.7605700, -1.2102626, 0.0115036, 0.5969367, 2.0109134, 0.3219413, 0.7599356, -0.2104610, -0.7714538, -1.9260959, 1.2535401, -0.0035488, 0.3836407, 1.0795503, -2.6641283, 1.7991973, 2.2081794, -2.0890227, -0.0457407, 1.2587249, 1.0986915, 2.3907571, -1.6297586, 1.2470508, -0.1607651, -0.1129111, 1.8697280, -0.2000908, 0.8203369, 1.8556651, 0.8959387, -0.1451558, 0.8585675, 0.4560811, 2.6095296, 1.2825918, -0.6396998, 1.7831431, 2.8456648, 0.7071261, -0.7282503, -0.0077861, 2.6222113, 1.1333045, 0.1394831, -2.2776735, -0.8938216, 1.5825066, -2.3736088, -2.7975086, 2.5650268, -2.7863443, -0.4571338, -1.1821026, -2.1547726, -2.9644958, -1.5884568, -2.4832503, -1.5886623, 0.3967865, -0.5886544, -1.4780107, 2.9319450, -1.6493285, 1.3486205, 0.6957411, -1.0684059, -1.0757850, -2.2666384, 2.4846739, -1.1868731, -1.2246808, -1.9217110, -2.6123458, -2.1595449, 2.1821883, 1.5386164, 1.1596580, 1.5666582, 2.5484619, -1.6128366, -2.5882454, 2.6396071, -1.6021851, -0.4791328, -0.6390679, -1.1781572, -2.1172160, 0.4296525, -0.6363686, 0.0624830, 1.7112260, -1.6712651, 0.9499575, -1.3793022, 1.7410440, -1.2482520, -0.0035399, -2.9916508, 1.5125191, 0.8779645, -1.8001397, -2.8773546, -0.1750491, 2.7335222, 1.9146766, 0.6960249, 1.0146091, -2.6634805, -2.9853356, 2.9395840, 1.9198806, 1.9992819, -2.4156951, 0.6383903, -2.3373076, 1.6883128, 2.1599018, 1.2062396, -1.0600678, 2.4131233, 1.9300503, -1.8717272, 2.8253330, -1.0610797, 1.3623000, 2.7443556, 2.9078587, 2.8375045, -1.6495332, -1.7134634, 1.1426720, 0.3293617, 0.4951223, 0.4974200, -1.9304372, 2.3918878, -1.7424640, -0.6292346, 2.7451349, -2.0686093, -0.9685437, 2.4885111, 0.9637206, 2.9055552, -1.6021883, 2.8765820, -2.7591224, -1.7732925, -1.8699947, 0.6626929, 2.5795833, -0.7388733, 2.0730925, -0.5096119, -1.6480824, -0.9528869, -2.6677604, 2.0009717, -0.4121233, -0.0480871, -1.8146929, 2.8807437, -1.6521883, -2.6862701, -1.5648432, -0.1888238, -2.3839651, -1.7275914, -0.4686272, -2.0134263, 2.8977071, -1.5841488, 0.1591044, 2.5543841, 2.9977793, -0.7770404, -2.6476183, 2.2021836, -1.6776779, -2.8071976, 1.8163091, 2.7648275, 1.4977237, 2.6876061, 1.9975935, -1.9289411, -0.8730930, 2.3781159, -2.5998961, -1.6912574, 2.7363117, 0.9849812, -0.7885166, -0.5382217, 1.0577737, 2.5967552, 0.2636381, 1.0410446, -1.6654305, -1.1462559, -2.6318504, 0.0562250, 0.8431237, -2.5224504, 0.2517177, -2.8853423, -0.0564646, -0.9508610, -1.2477502, 1.1978336, 2.9623023, -2.2140833, 1.9516587, -2.5468868, 2.8286996, -1.2474364, -2.3271027, -0.9394422, -2.4110709, -1.7674685, -0.0401922, -1.6571056, -1.3107237, -0.9656139, -2.4270385, -1.4704042, 2.5938015, -0.6470534, -1.3044415, -2.5781720, 2.8451612, 1.1340723, 2.4886130, 0.7400633, 1.3440546, -1.2834696, 1.9717252, 1.2427618, 2.6386699, -2.9362162, -1.1019387, 2.9780741, 0.1725828, -0.4151827, 2.4747795, -2.1467722, 2.1228542, 1.1226205, 1.8241688, -0.9071568, -0.0109673, -1.3768710, -1.1675744, 0.4738936, 1.2118783, 1.6705476, -0.0306596, 1.0766024, 2.6522629, -0.1534189, -2.7078974, 2.5333520, 1.5085999, 2.3097271, -1.1797895, 2.4672319, 0.8971363, 2.9204611, 1.0955871, -2.3653802, 2.3059669, 1.1021749, 0.4097272, -2.2365987, -2.2232416, 2.1110526, -1.7581428, 1.1801450, -0.5329242, 1.9166199, 1.0637141, 1.5892418, 0.3228033, -1.3914311, 2.8695006, 2.2615654, -1.4986130, -0.2309509, 1.1242825, -0.6065650, -1.3096029, -2.0834335, -2.8568100, 0.3849390, 1.1751749, 1.8972011, 0.9138762, -1.5575662, 0.5330724, 2.8544866, 1.4100299, 2.1509749, 2.2901674, -2.8468257, 2.0926803, -2.0516347, 2.6880803, -2.7093320, -2.3742996, -2.9323345, -2.7156591, 0.3316689, -0.7981818, -2.7103964, -0.6788924, -1.2350110, 2.7076333, 2.0141612, -0.1769067, -0.7183203, 0.3337307, 0.4071996, 2.9656582, 1.3436574, 1.7454868, -1.8093288, -0.2514504, 2.8856017, 0.6646247, -0.2520726, -1.4176662, 2.5519366, 2.8223697, -2.7676988, -2.0522158, 0.4923120, 2.8769451, 2.4740554, -0.2918816, -0.4132585, -2.3582541, -1.5323205, 0.8841032, -1.7578599, 1.8959394, 2.3836288, -2.2785352, -0.2769730, -0.7267666, 1.3866864, 2.3440105, 1.9128248, 1.8877528, 1.4864434, -2.2148052, -0.8374083, 2.2529159, 1.6502616, 1.9287579, 0.9622425, 1.4482791, 1.1543095, 2.1685545, 2.2259724, -1.4611967, 0.2591029, 1.1614151, -2.8081532, 1.5611877, -0.3124218, -2.3742182, -2.9277859, -1.3474925, 0.9914956, -2.2319284, 1.1085464, -2.1122544, 1.1110085, -1.3646882, 0.2428232, -2.3852357, -1.6189029, -2.5836503, 1.7120074, -0.3548492, -2.1202841, -2.4580711, -2.4967145, -0.3044599, 2.0264229, -1.4919094, 2.6532242, -2.7774581, -1.8280442, 1.9686464, 1.6338943, -1.4560796, 2.3353697, -1.8384831, -1.3169512, 2.7201561, 2.3901547, 2.0495597, 1.7899582, -1.2073478, 1.4361572, -0.0829983, 1.0464117, -2.3457453, 2.3146016, -0.4076858, 2.5392910, -1.7903586, 0.9080995, 2.2669837, -1.2160239, 2.7273284, 1.8232701, -1.2905765, 1.0493512, -0.0281857, -0.1520517, -0.1410572, -1.9528176, 1.8608466, 1.6162127, 2.7433807, 1.3294788, -0.1242168, -0.6633441, 0.0511691, 2.6580583, -1.7917972, -0.7728150, -1.3197936, -1.5604541, 2.2546938, 1.0661404, -0.6972972, -0.1720178, 2.3173847, 0.2335158, 2.9900759, -1.3940115, -2.3492612, 0.1686802, -1.5193399, -2.5028299, 2.1238806, -2.8510527, -0.7271157, 2.1867106, -1.8996811, 0.8827260, -0.2024843, -0.5005702, -2.5358053, 1.9535621, 1.0716941, 2.8922303, -1.4769504, -2.7915161, -0.7722811, -0.8802693, -2.6149148, -0.2761081, -2.2931985, 2.7625587, -2.5699877, -2.6841790, -0.3266997, -1.5577098, 2.4860786, 0.2778983, -1.7076187, -1.3843838, -0.7991376, 2.4158763, 0.7352595, 2.7514510, -1.8594089, 1.0767976, 1.9969362, -1.8078183, -2.8630604, -0.0184519, -0.4433034, 1.8934424, -0.2959976, -1.5538795, -2.1730788, -0.4141317, -0.8099436, -0.7884599, -1.3785402, 1.7271026, 2.9816646, -0.1883411, 2.9430948, 1.9334006, -1.3711884, -0.7297858, 1.7792136, 1.2343450, 1.0215568, 2.7482941, 0.1199445, -0.1104580, 2.8925433, 2.3437197, -0.5332621, -0.1899110, -2.0986702, -1.1636142, 2.3388237, -1.7269913, -2.3181499, 1.4510646, 1.1479540, 1.2435438, 1.9292381, -1.7098209, 1.0105675, -2.6585747, -2.7169844, 0.4640120, 1.4322766, -1.6590266, 2.0268967, 2.2421918, 0.1054433, 1.5398956, 0.5919515, 0.4990058, -2.8669190, 0.3625844, 2.7244739, 0.6554675, -1.2662251, -2.5149767, -0.4078734, 1.2302839, -1.5740359, 0.3183531, -2.7716975, -2.7640897, 2.2931951, 2.6817732, 0.1180011, -1.2942545, 2.1456801, 0.8160053, 1.1873767, -2.9294490, -2.7381541, 0.1371545, -1.3113955, -2.0599468, -2.7513170, 1.5253305, -0.5500360, 1.2662383, 2.3194350, -1.9554819, 1.7598349, 0.1066743, 1.8482834, 2.9946768, -2.8893921, 2.3222131, -1.4719459, -0.4861319, 0.5139886, -2.0851013, 2.1396391, 2.6045805, 0.9238745, 1.7830696, 1.5812403, 1.1343729, 0.9197133, 2.5629734, 1.2181324, -1.7909953, -1.5943816, -0.8862621, -0.3567475, 2.3098680, -1.3297334, 1.5973952, 0.3810182, -2.0114307, 2.0831091, 1.0836294, 0.3243100, -1.2648211, 1.6769994, 0.2178850, -1.8608640, 2.8599423, -1.3999684, 1.8025237, 2.3041580, -0.3298072, 0.1198610, -2.1895693, -2.2060549, 2.6246987, -2.8395391, 2.3343271, -0.0686519, 2.5677601, -0.5297255, -2.4244149, 2.5553546, -1.0513735, 0.8001812, -0.2407724, 2.4981278, -2.7745824, 0.9222646, -0.4233826, 0.0231621, -2.0928161, 1.4108375, -0.6971399, 1.5967466, 1.4787889, -2.7993111, 0.7252980, 0.1588863, 1.3801216, -1.2640894, 1.7090900, -1.8030457, -2.7726044, 0.1931468, 2.6262423, 0.3789628, -2.5512953, -0.6783607, 2.3332565, 0.5263400, -0.6347556, -0.6995819, 0.6290438, -0.2827733, -0.6298781, -2.7272756, -2.5293701, 0.4635073, 0.2930711, -2.7872809, 2.7566656, 2.7003101, -1.5741236, -0.9637208, 1.2124762, -0.8924081, 0.5363262, -0.9260962, -2.6470911, -0.7827207, 1.3290247, 1.4239558, 0.6237641, 2.4609468, -0.8038041, 0.8145908, 1.3347575, -1.4726482, 0.5265280, -2.2885998, 1.4222271, -0.3956209, -0.3064219, 2.7728827, -2.5322755, 0.1469662, -2.3567342, -2.0271694, 1.9942951, -1.3533627, -1.5600144, 2.0857004, 1.8207972, 2.7283114, -1.9089184, 2.5196264, 1.3772880, 2.6556700, -2.3905635, -1.3571562, -2.0437421, 1.4553339, 2.2515355, 0.7964857, -0.8471592, 2.1752911, -1.0783284, -2.6010547, 2.5816295, -0.9493635, 2.9917046, 2.8560009, -0.7611494, 2.8923852, 1.9623440, -2.1265511, 0.2189827, -1.1054105, -1.3883576, -1.2139229, 1.2922676, -1.0087256, 0.5048549, -1.5277515, -2.3322964, -2.5718100, -1.5807429, 0.4454739, -1.9222117, 0.9244708, 0.1081290, 1.5989239, 0.3116547, 0.4896602, -2.8627708, 0.3255834, 0.4311920, 2.1960873, 2.7073385, -0.8610266, 1.6834574, -2.5841564, 1.1770361, -1.7877572, 2.7044392, -2.1080460, -1.3871376, 0.0171507, 2.2314112, -0.0099101, -2.4696486, -1.6734320, -0.8154998, 0.7197729, 0.3677269, -0.9523685, 1.2121700, 2.6358939, -2.7736000, -1.0204686, -2.2699671, 2.7490588, 1.5784215, 0.9220732, 1.7449226, 0.7542777, 1.3414112, -0.4001740, 2.9397266, -2.1836849, 2.2819744, -0.3723596, 2.3514931, 2.7727087, -0.7185430, -0.7258846, -0.8589393, -0.0724804, -1.9916795, -1.0329208, 0.2746018, 1.1418404, 0.7254480, -0.0997060, 2.6723271, -0.6386976, -1.9287385, -1.6732046, 0.3131858, -1.2132532, 0.0568361, -0.5238235, 1.0694808, -1.8583639, 0.2368674, 1.5837507, -0.2548848, -1.1451051, -2.3394063, 2.3518701, -0.9106596, 0.3749219, 0.4764155, -2.9589324, -0.9865924, -0.6546910, -2.4666146, 1.9457465, -1.3145872, 0.4331390, 2.9872346, 0.7615640, -0.1321663, 1.7611353, 0.7250453, -2.5732398, -2.5027544, -0.2073150, -2.2256399, 0.6901877, 0.8753012, 2.2807719, -2.3859548, -1.9622083, 0.0491427, -0.4550357, 0.4824086, -0.4773962, -1.8972324, 0.5497605, 1.6323894, 0.4656774, 2.3209369, 2.1184986, -2.8670322, -1.3720861, 0.8224909, 2.7694085, 1.6224737, -2.2171891, -2.3765774, 0.4614840, 0.6915900, -0.7267927, 1.7345280, -2.7032516, 0.9698162, 0.4380506, 1.9883091, 2.5022433, 2.9076406, -0.5450641, -0.9920158, 1.2603046, 2.4993952, -1.9615778, 2.8964662, 0.8656034, -0.3357039, 2.5094338, 2.0553608, 0.1456869, 0.1069924, 2.8673398, 2.3075694, 0.5981155, -0.6179752, -2.4804915, -0.0970757, -1.4407677, -2.6520821, -2.5408818, -0.1440399, -0.1944941, -2.4254870, 0.0952908, 0.2817307, -0.5656970, -0.2048231, -2.3093090, -2.5144645, 2.2433201, -0.7453534, -0.0780003, -0.7904040, 1.5249669, -1.7964088, -0.7794956, -0.4395900, -1.7588387, -0.6239793, -2.6953636, -1.5748761, -0.9166330, -1.1518965, 2.4520743, -1.9941729, 1.7374836, 2.0053262, -2.1169605, -2.1785911, 0.7153500, -1.0600041, -1.7490511, -0.3557863, 0.8983251, 1.3138343, -0.7489557, 2.9739466, 2.0482689, -2.5171478, 0.9071530, 2.9547687, 1.7274299, -1.9571365, 1.7130966, -1.1790205, -1.4094581, 1.2678124, 1.0946524, -2.8262611, 0.1010629, 2.6293994, -2.5318069, -2.1094196, 2.1011858, -1.0716156, 0.2154277, 0.7919120, -1.6496380, 1.8787502, -2.8960551, -2.3206101, 1.6546281, 0.8649980, -2.4153330, -0.7486343, 0.9009053, -2.5915534, -0.4943941, 2.6561874, -0.7878037, -2.0282770, -1.1310712, -0.6206580, -0.7253789, -2.4814652, 2.9781255, -0.0620366, 0.4997458, -0.4960608, 1.0101991, -2.1250440, -2.8182832, -1.8927876, -0.3375732, 0.7195705, -0.7372752, -1.0647446, -1.7681088, 0.6402654, 2.2564512, -2.5545049, 0.6872017, -1.9880109, -0.6620968, -2.5717650, -0.4456596, 2.3188349, -0.9919097, 2.3189775, 2.0297487, -0.7367743, -1.6063068, 1.1334205, -2.1107585, -2.8788270, 0.6188119, -0.1343680, 0.0084425, 1.7433591, -0.2596723, 2.4111049, -1.8986542, -2.6283116, -1.0842415, -0.5080558, 1.4278398, 0.0823983, 0.9000119, -1.4501480, 1.6196263, -1.7542400, -2.2469100, -1.3889783, -2.0414847, 2.7084152, 2.7271422, 1.1425280, 2.2950176, 2.1912774, -0.2470347, -0.4749195, 0.5323139, -0.3928519, 1.2365723, 0.3980505, -0.6985425, -1.9623680, -0.3275384, -2.8609700, -1.6838776, 0.2825726, -1.8124770, -1.3512285, 1.1047098, 2.2589395, -2.8268083, 0.1589006, -2.6082201, -2.1487461, 2.9248556, -2.2671427, 0.6884207, -2.9098577, 0.1403309, -2.3810586, 1.0418955, -2.7413230, -1.5516085, -0.4762787, 1.6169639, -2.6854537, -0.0746028, 2.8145243, 0.5417811, -1.9964471, 1.8979767, 2.9004446, 1.0695585, -0.5547128, -0.3992470, -2.7283460, 2.1825937, 2.6229478, -1.3433577, -1.3276068, 2.8280835, -1.2505454, 1.3724308, -1.6590797, 2.1115311, 1.6435302, 2.2891745, 2.4798789, -1.8802651, -2.2410574, 2.8370629, 2.2655109, 0.0057182, 2.4700084, -0.4537528, -0.5912363, -0.4944665, 1.1318038, -1.3533395, 0.4498702, 0.0877774, 0.3220638, 2.3417927, 2.8414848, 2.0243694, 2.0275498, 1.6434416, 1.8197313, -2.7298649, -1.8396209, 1.8885668, 1.0429499, 2.2502097, 1.6907560, 1.7578307, -0.3241569, -2.7410085, -0.8400816, 1.1743811, 2.8047625, -0.3606361, -0.6461308, -0.2543624, -2.6370504, 0.5552503, -0.7208776, -2.9115492, 2.2110486, 0.4363002, 0.1682136, 1.8025548, -0.6595794, -0.7745559, 1.1702830, -0.0121658, 0.5676020, -0.5833525, -2.5008248, 2.1260643, 2.7132364, -1.5299628, -0.2870781, -2.0402680, -1.5558138, -1.8449869, -1.7032524, -0.7715796, -2.5104062, -2.9799955, 1.1239569, 1.3621510, 1.7378987, 2.7992269, -0.7169322, -0.3767147, -2.0733621, 1.6021596, 1.4925268, -1.0447890, 1.1017832, -2.4615748, 1.2928503, 1.2142837, -0.8700227, -2.5250944, 2.0415992, -2.3351987, 1.9361638, 2.2746983, -1.9051055, -2.6696856, 2.7052004, -1.9941610, 0.0057582, -0.6221470, 0.9849172, -2.9049069, 0.0947859, -0.8246899, -0.1245070, 2.7039008, 1.6637495, 1.9962968, -0.2298933, 0.2693169, -1.0422400, -2.3767314, -0.3180390, 2.6761863, 0.6711872, 0.2934473, 2.1291866, -2.8645401, -2.1102490, -1.9349563, -0.0503350, -0.9632954, -0.0520629, -1.1556241, 1.6323281, -1.6841576, -2.5791948, 2.1881398, 0.8609751, 1.0325579, 1.3111816, -1.0880510, -2.3848016, -0.3243392, 0.5766134, 2.3920912, 2.2531352, -0.4095048, 2.1990130, -0.0056300, -1.5301838, -2.7481028, -1.8868367, -0.0369903, -2.9436620, 2.4554065, 2.4025642, 0.6529968, 0.2407018, -1.5540892, -2.6976760, -1.7614000, -2.2080071, -0.3336932, 1.2260102, 1.5629699, 1.1168174, 0.9175992, 0.5963026, 0.1798671, -1.2907586, -1.8855488, 0.0638955, -2.9575297, -1.4200479, -1.6433107, 1.6858530, -1.1344261, -0.6225512, -1.9998171, -0.0949195, -2.6745244, 1.5654482, 0.3394212, -1.3608278, 0.8834263, -1.8053976, -0.2212253, 1.4345265, -0.3209509, 2.7121971, 2.0409035, 1.6871308, 1.4276766, -0.1417160, 0.3511196, 2.1235724, 0.1716303, -1.6580814, -2.6807318, -0.5029004, -2.1260271, 0.4511235, -0.6436225, -1.5075011, 1.8734935, 0.7296567, 2.0248200, 0.8922823, 2.5865143, -0.4462095, -1.2551947, 1.3478191, 1.2784291, -1.4376028, -2.8268515, -0.8853952, -0.0961953, -1.3919055, -0.9839727, -2.5607210, 2.7107986, 1.0647625, -1.7359190, 2.4197697, -2.6610249, -0.5873878, 2.7993404, -0.5878002, 1.1047890, 0.9168608, -1.7015242, 1.2580579, 2.1342715, 1.3666102, 2.9425520, 2.3208457, -1.9376507, -0.3829767, -1.1549691, 0.7381680, 0.3957312, 2.7902333, -2.6946634, 0.4492589, 1.4034684, 2.8495927, 2.8119971, -2.2570528, 1.7727721, -2.5616038, 1.5728367, 1.4969279, -0.3408040, 0.2437148, 1.8454583, -0.5561602, -2.7200252, -0.9644899, -1.7066925, 2.6184299, -1.9194084, 1.2659946, -0.6591202, 1.4278803, 1.4822164, -1.1586604, 1.9823772, 2.4612078, -0.3175097, -1.2474003, 0.1023009, -0.0678682, 0.1195103, 1.9389580, -2.3401923, -1.8777633, -0.9058682, -2.6404641, -2.6167743, -0.0366665, -0.7524458, -1.0350305, -1.6853516, -2.7036536, -1.2797865, 0.2424391, -0.3561221, 0.6162021, -1.4990817, 0.8051859, 0.1883628, 2.6464814, -2.6702467, 2.0294821, -0.2599083, -0.6823749, 2.7812854, 2.7475400, 2.4342225, 1.8096831, -2.2526563, 1.8912545, 0.4162666, 1.1741523, 2.7435121, 2.9862600, -0.9789227, 0.7145061, -0.0997342, 1.1880373, -2.2838158, -0.5220126, 0.1751576, 2.2526946, 1.2574315, 2.9155717, -0.8843915, 1.9534551, 1.5412764, -0.0403627, -0.7306102, 0.3852783, -0.3985337, -2.5869049, 2.7145463, -2.5800991, 1.5786727, -2.3979052, -0.5945751, 0.7176213, -0.9784380, -2.4931488, -1.7003281, -2.2655344, 2.4692571, 0.7917647, -0.6533513, -1.6269178, -1.5451263, 0.1936968, -2.9985399, 1.2836572, 2.1623602, 2.2409631, -2.2007133, 0.3648624, -1.0611070, 2.2358635, 0.2717038, -2.9497772, -2.0262003, 1.8572572, -1.6592621, -1.0201947, -2.9835207, -0.1072191, 1.5895812, 0.5437574, -2.2177549, 1.5574700, 1.6370279, -0.9120259, 0.9772348, 1.6256183, 0.5885113, -0.2008039, -2.2238932, -1.4355227, -0.9407502, 2.3211888, 1.4781333, 2.9171398, 2.5627070, -1.4264177, -2.1652179, -0.2430347, 0.5622471, 1.5340882, -0.5310216, 2.2236797, 0.1476085, -2.5631407, 1.1968031, 0.4536981, 2.7857906, -1.3884320, -1.7827516, -1.3568503, 2.6643517, 2.5699212, 1.2055298, 2.0287238, 0.8901875, 1.4725204, 1.9232358, -0.8340420, 2.1186181, -1.9648178, 1.7647403, 2.0887367, -0.4150364, -1.0825662, -0.1020176, -0.1204294, 0.7120492, -1.3954016, 0.5737465, -1.2779251, 2.4638691, 2.6696849, 0.1086416, -0.6266861, 2.0202597, -2.9304471, -0.4160314, -2.9356674, 0.3722053, -0.4114810, 2.5620316, 2.4220022, -2.5892930, -1.5716139, 1.4449218, 0.8933324, -1.9276555, 0.5169706, -0.2163999, 0.2698412, 1.8918070, 0.0162358, -0.8256818, 2.7094289, 0.0260954, -2.0120440, 1.0049926, 1.6144157, -0.2173457, 2.8969767, -0.5639367, 1.9241903, 1.0736771, -1.7405876, -0.3037792, 2.2199080, -2.2799445, 2.7150277, 0.3239105, -0.9129050, -0.1852834, -0.5624722, 1.7269173, 0.2563646, 0.9196633, 2.7191294, 1.9715160, 0.9111079, 0.1009878, -1.6127893, -2.9744108, 2.3839502, 2.6795980, -2.6305340, -0.8435205, 2.2961129, -1.9884253, 0.9607742, -0.1894946, -2.0865309, -2.4019058, -0.4068291, -2.0191055, 0.7330868, 0.7154200, -0.6727790, 1.2811197, -1.7147856, 0.4813464, -1.1597127, 1.7110854, -2.7229877, 0.7411219, 1.2044512, 0.7513764, -1.9163407, -0.6537578, 0.2934949, -2.7509201, 0.7176251, -0.1958695, 0.7790260, -0.4843122, -2.8472863, -0.0649157, 0.0208902, -2.7366274, 1.4432445, -0.8263652, -0.7457332, 2.4385151, -0.7603392, 0.0525597, 0.3128819, -2.1322007, -0.1594114, 0.5502657, 0.0455073, 2.3250612, -0.8105447, 2.7602849, 2.7534423, 1.6756181, 1.5965751, -1.7843884, -0.6355361, 2.8580420, 2.4036032, -0.2410819, -2.6299609, -1.4180026, 2.9597676, 2.5732910, 2.2497897, 1.4378736, -0.5402754, -2.4694699, 2.1949962, 0.4301105, -0.8363638, 1.0704583, -0.2292273, 2.5306211, -0.6790208, 0.2602387, 2.8193006, 1.0669303, 0.3556117, -1.5936806, -2.3770589, 2.0720247, 0.2821742, -1.2130344, -0.1157540, 2.2430382, 2.1216748, -2.5624729, -2.0000108, -2.5376806, 1.0445494, 2.1477133, -1.1335045, -0.4437736, 1.1217102, 0.7467411, 2.7532997, -2.5025652, -0.7695790, 0.1536531, -2.3660802, 1.3088806, 0.3978842, 0.9333559, 2.2428666, 0.5237028, -2.7278533, 2.4251363, 1.5605231, -2.4614968, -2.4509237, 0.3634325, -0.8134148, -1.4119128, 0.1031219, 2.0784453, -1.1186266, -1.7465892, -1.5441477, 2.1453125, -1.9013890, 0.5215239, -1.7930315, 0.0577716, 0.1666611, -2.0226311, -2.1460949, -0.1083645, 2.4854718, 1.5248473, -0.3208019, 2.9542333, -1.6452841, 0.8634022, 0.7849436, 0.4030592, 1.9321800, -1.7786125, 2.7546733, -2.5063654, 1.1353161, -1.0177114, -2.8540931, -2.9643353, -1.2608962, 1.6676601, -2.2861188, 0.1421495, 2.1486427, -2.4570649, -1.8276338, -0.9239498, -1.4238283, 1.8962289, 2.6930085, 2.4637814, 1.2134779, -0.8891608, 0.5187751, -2.7879785, -2.5199752, 0.2921681, 2.3387040, 0.2314887, -0.3325871, -2.9218177, -0.8829570, -1.1218969, -0.0779216, 2.6166080, -2.7886644, 0.0963782, 1.2600901, -0.8165772, 0.5845396, -1.4631535, -2.0404264, 2.1542742, -1.3344035, 2.1958617, 2.9337597, -0.8943471, 0.1592971, 0.1731544, -0.4316520, -1.6254913, -2.5943079, -2.1253535, -1.3954392, 1.5655382, -2.8571005, -1.7270466, -2.5297114, 0.4074862, 2.7810311, -2.5351826, 1.6399361, -1.3467362, 2.2586501, -0.7485344, -1.5896333, 1.4562155, 0.4573284, 1.9494848, 2.5765766, -2.9442430, 0.5059540, 2.5893164, -1.7260973, 2.8940747, -1.1997291, -2.2145594, -2.7619905, -1.4406926, -1.9366400, -0.0000463, 1.5097801, 0.6750873, 2.8360855, -2.8242145, -2.0402745, -0.4883474, -2.0098819, -0.5538933, -0.4883665, 0.0883389, -2.6555789, -2.0479502, 0.9502314, -1.7144237, 0.1522209, -1.2543877, -1.9945686, -1.8191773, -2.9732597, 1.4404277, -2.6162201, 0.2027397, -1.3536679, 0.8478753, 2.9251910, 2.6582589, -2.7224479, 0.8868822, -1.0882507, -2.4834311, -2.5457902, 0.5783422, -1.2625238, 2.4254506, 1.4806853, 0.6817048, 0.4828091, -1.4971421, -1.7681418, -2.1649658, -2.3465257, 1.3002216, 2.1083827, 2.4350315, -0.9784681, 0.8019094, 1.9070086, -0.1641762, 2.5451660, 2.0609599, 2.5915151, 1.0949454, 2.4352013, 1.7362275, 2.4620028, -2.3200681, 2.9337197, 2.8738975, -0.6582226, -0.2013837, 0.1403482, 1.5086811, -0.4900091, -0.0218109, -2.4755453, 2.5965481, 0.6572953, -2.6560469, 0.7410847, -0.6878265, -2.7949149, 2.7774470, -0.8154626, 0.3235073, -1.0845980, -1.2544783, -1.8456410, -1.0056965, 2.9685437, 1.4431367, 1.1362126, -0.3260228, 2.7973388, 2.1635347, -0.3607408, -1.2368534, -2.1059467, -1.4058388, -0.8187294, 1.1987283, -0.9364989, 1.8003998, 0.4809103, -2.3638050, 1.6905065, -2.6062644, 0.3616986, 0.6124515, -1.9503602, -1.0739502, -2.4824661, -2.9652988, 0.5706637, -1.2479729, 1.4776442, -1.3664069, -1.6116017, 0.8522483, -1.5151424, 0.7697356, -0.0906263, 0.5607903, -0.2245268, 2.8108639, -1.9531920, 2.6055207, 0.9025580, -0.3308603, 2.5585331, 1.5903883, 0.1759780, 2.0074661, 0.6155549, 0.2001512, -1.3867640, 0.5768787, 2.0301336, 0.1312094, -2.7166759, -1.8378480, 1.9563014, 2.3738043, -2.6633280, 2.6418645, -2.1929487, 0.9267580, 0.5862241, 0.7305414, -2.3033741, -1.4001511, 2.7926084, 0.5392804, -1.7928152, -0.5455565, 1.6802393, -1.6318055, 0.8189471, -1.2312063, 2.8214663, -1.1510279, 2.6559163, -0.4509338, -0.2480775, 1.4439097, -2.1353622, -0.0800106, 1.3038036, 1.0705967, -2.3796167, -2.6985612, -0.1790635, -0.4621205, 1.3899570, 2.6084474, 2.2431768, -0.2154300, 0.6720056, -1.7747365, 1.4426936, 0.6871688, 2.4807965, 2.1525670, 0.0964088, 1.7962600, -2.2956702, 0.6840113, -2.1762841, 2.3104488, 0.8979974, -1.2045055, -0.8561962, 2.0463625, 2.5524978, -1.2797777, -0.3710956, 2.7085954, -0.6382078, 2.5321470, 2.0377836, -0.5463874, -2.4566112, 1.0164974, -2.3827668, 1.3941800, 0.2318006, 2.7672966, -2.4601833, 0.1007672, 1.1687037, -1.2099124, -1.8271168, 0.4671861, -2.3650871, 0.4001004, -1.3236737, 0.4938633, -0.5814219, -2.2721082, -0.3551780, 2.1910104, -1.1061454, 2.5858627, 1.3321365, 0.1844984, -1.6629164, 0.6571207, 2.2649013, 2.4264832, -2.0524121, -0.9931697, 2.1608971, -0.1653077, 0.1849534, -1.2037769, -0.1417997, 2.9280358, -2.9937445, -1.5411619, -1.8408243, -2.6849842, -2.8796514, -2.0485388, 1.8245125, -2.5163442, -0.3624793, 2.3934203, 1.3461188, -2.1707557, 0.0014289, 2.4356591, 0.1597001, -0.9510611, -1.7359067, 2.1137281, -2.3665319, -0.5239197, 0.2618727, -0.5344625, -0.1583612, 1.4718260, -0.2220502, 0.1802932, 0.8740239, -2.2045053, -2.7277274, -1.9818335, -1.1190597, 0.7942937, -0.1381265, 2.8533185, 0.6928533, -2.2709054, 1.1405677, 0.5738138, 2.0423060, -1.8078415, 2.7481730, 1.6494053, -0.7844260, 0.3377533, 1.2945919, -0.9211093, -1.5539744, 1.5691980, -0.4791106, -1.9548415, -1.7094863, -2.7464533, -0.2324540, 2.3012214, 2.5917679, 1.6345341, -1.9993867, 0.8512834, 0.4738685, -2.9574990, -1.3450529, -0.7057859, 0.2100705, 0.8679986, 0.9177757, 1.8138420, -1.6399633, -1.8253496, 1.4120639, 2.1674288, -2.9930662, 0.4800378, -2.7815612, -1.8602037, 2.9469324, 2.8809771, -0.9853103, -2.0763591, -0.9993730, -2.7924347, -0.3541909, -1.2940034, -2.5802796, 2.4770373, 0.3704440, 0.9651808, -1.7933984, 2.4771942, 0.3209480, 0.1427556, 2.8220494, 1.9352694, -2.1901184, 2.0120268, 2.5946097, -1.3330035, -0.7099424, 0.5031359, -1.1988894, 1.0450410, -2.3941222, -2.9427733, 2.1173703, 0.2422800, 1.2356781, -2.3394224, 1.3938038, -0.9987983, -0.3417272, 2.1432365, -0.8325539, -0.8602559, 2.1106999, -1.6170871, 2.5442977, 1.4103559, -2.9787267, 2.1748479, 2.6936459, -1.1976716, -0.5778280, 2.3932418, 1.1455116, 1.9820674, 0.4398971, 0.3470492, -1.7533257, -1.5451925, 0.9965871, 0.9322867, 0.0869096, 0.7444812, 1.9013252, 0.5066505, 1.6136857, 2.2876281, -1.3968084, 0.7039542, 2.5888234, 1.5450737, 0.5253430, -2.7733677, 2.7356150, -2.3426490, 1.3793942, -1.5971842, -1.1616167, 2.1434273, 1.8771956, -2.1040923, -1.7929337, 2.9356120, 0.6826957, -1.0829041, 0.6674275, -0.9069742, 2.8560722, -0.0024370, 2.2620044, -1.3143049, -1.1297103, 1.0871422, -2.8729783, 2.8862985, 0.8505853, 2.5120615, -2.6650952, -0.2883019, -0.8920652, 1.1216158, 1.2309069, -1.3534763, 2.3045436, -0.8123336, 2.0173053, 1.3661283, 2.3183343, 2.1662609, -2.1453836, 1.5674906, 1.7509874, 1.4943867, -1.8006187, 1.9111506, -0.6966039, -0.6167136, -0.0902441, -2.1893474, -2.6778271, 0.2226105, -2.4212795, 0.7425441, -2.2441326, -2.9455895, 0.8930342, -0.2410320, -1.2064432, -2.4795466, -2.3457348, -1.7946991, -1.3636146, 2.0739275, 2.4541504, -1.8156437, 2.6074851, -2.3200573, -0.4086035, -2.2719433, 2.8327747, -1.7265044, 0.2545642, -0.9544900, -2.2425059, -2.8812723, 1.0476112, -0.8401309, 0.0363831, -1.2953874, -2.6525673, -2.2463031, -2.1108360, -2.4017453, 0.5953544, -0.2313056, -2.2304506, 2.8901553, 2.0770425, -2.3396872, -0.2987595, 0.3196915, -0.4738368, -0.2956321, 0.2109985, -2.7817606, -0.2661662, -2.4658687, 0.4288492, 0.5510696, -2.5268300, 1.3451342, -2.7122102, -2.4913985, -1.6086175, -0.4451802, 2.0857135, -1.4456752, 2.1461153, 0.7859517, -0.3182348, 2.6603806, -1.6965311, 2.9813728, -2.5363796, -0.8720759, -1.1063043, -0.7557075, 2.7113376, -2.1368245, -1.8457855, 0.0240706, 0.2874654, -1.8646358, 1.2339299, -1.5656736, 0.1478682, -2.6018907, -2.4076642, 2.4509768, 1.5756317, 2.8203192, 2.5703436, 0.5762988, -0.0218209, 1.6178310, 0.3822085, 0.5167456, -2.6161223, 2.7916027, -1.8656020, -1.9323002, -1.5147556, -0.0303801, 2.0191680, 2.4775183, 0.0948439, 2.4188864, -2.9361967, 0.0958726, -1.7180265, 0.9988516, 1.0481378, 0.6234059, 2.8536867, 1.3951058, 1.8861386, 0.8122613, -1.6007087, -1.4348046, -0.0417432, 0.3773232, -2.9348146, -2.6083989, -1.2270734, 1.1791206, 0.4045612, 2.7204762, 1.2831622, 2.7765673, -1.4701495, 0.7185052, -2.2991713, -0.3330033, 0.7767811, 2.3744110, -1.0236936, 0.5785138, -1.8947359, -0.5324212, -1.2551833, 1.7294229, 1.9129727, -2.9652501, 0.1896992, 1.6216978, 2.7889369, -2.6982837, -0.5645958, 0.8684002, 1.5048387, -1.6378242, 0.6433236, 1.4878831, 0.9533548, -0.7107923, 2.7898998, -0.9933901, -1.5630123, 1.4544721, 2.6685789, 2.4044950, 0.6571448, 2.2691208, -1.1572081, 2.8312529, 1.2010991, -2.1335685, 0.5695718, -0.5533980, -2.7642933, -0.4013353, 2.8436002, 0.1355043, 2.1425481, -1.2430454, -1.3886425, -1.7198742, 2.2822978, 0.9425187, -2.5500863, 2.2062512, -1.1084781, -0.6644008, 0.2850199, 0.0651582, 0.9045959, 0.3407200, 0.1194874, -0.3385977, -2.4746506, -1.7578749, -2.6977036, 0.4170048, 1.3363832, -1.2042169, 2.3128742, 1.9601586, -1.2997359, 1.9021484, 2.8091260, 1.5353429, 1.1774773, 1.6803588, 0.0826702, 1.1877330, 1.3628664, -0.3262326, -0.0393575, -1.0054726, 0.9399903, -1.3894793, 1.2953195, -1.7398494, 2.9086526, 0.6836035, 1.5169537, -2.4249369, -2.3457644, -1.2807011, -2.7165967, -1.9717887, 1.7075360, 1.5678138, 0.0305058, -0.7336817, 0.4960183, -2.8150598, 2.8080639, 2.8207683, 0.1961135, 0.3943704, -2.7916606, 0.7511853, 2.3332246, 0.2664671, 1.0978729, -0.8069987, -0.0230527, 0.9093693, 0.1550058, 0.4075007, -2.7371044, 0.9662926, 0.4549836, 1.9010892, -1.7447916, 0.9133728, 2.3704065, -0.5182394, 1.8067737, 1.2776992, -0.6476364, -2.2021753, 0.0174995, -1.3585409, -2.9376920, 0.7556708, 1.4819554, 0.7222590, -0.9759451, -0.1606033, 0.0422737, 1.1608511, -0.7196120, -0.9212562, -1.5368194, -0.1876898, -1.9347478, -2.6782362, -1.5507059, 0.4747207, 0.3505766, -0.1523726, 1.0455594, -2.1250845, -1.1013560, 0.7522311, -0.7736163, -1.8673263, -0.6764144, -2.1607017, 2.4086469, 0.8216300, -0.7424793, 1.1961487, -2.7080723, -2.1369786, -2.1558295, -2.7497909, -0.9808434, 2.2085726, -1.2671344, -2.2890520, -2.1014864, 1.0522780, 1.8449879, 2.3993801, 2.9597940, -2.9401399, -1.5497816, 0.6568523, -1.2448307, 0.5348702, 0.9499796, -0.9169778, -1.5577753, -2.9121705, -2.6470856, 2.9769383, 2.2782783, -1.8099182, -1.6585228, -1.0509000, -0.6894569, -0.8601329, 1.5153364, -2.7021764, -2.4577796, 1.3925061, -0.4023956, -2.1051040, 2.2081796, -1.6363495, -1.9718801, -2.1155334, -0.7028128, 0.2669341, 1.5892598, -1.2413839, 2.0133166, 1.9593721, 2.9855198, -1.8610433, 1.5833759, -0.9396555, 2.1753132, -1.1761006, 1.1485175, -2.2352069, 1.5327696, -1.9000392, 1.5785575, 1.2731875, -0.3310094, -2.4717255, -1.3143000, -2.9461782, -0.8803269, -1.5003050, -1.7929636, 2.0112716, -0.2444869, 1.9714176, -0.3736031, 0.7584748, -1.7791544, 0.4988459, -0.7671012, 1.4644488, 2.1972283, -1.0848738, -0.9331935, 0.8366621, 0.6083628, 2.5692507, -2.7506654, -2.6145236, 2.3347840, 0.4425383, -2.1548129, 2.3804471, 2.7963655, 1.0534215, 0.5084349, -1.7035561, 0.3644531, 1.7609341, 2.1557289, -1.7649545, -2.5352441, 1.6033353, 2.8052666, 2.3437641, 1.6762651, -2.3135178, 2.8878185, -0.7016790, -2.1488667, -0.3337517, -0.4591118, -1.0994202, 1.2379876, -2.2472293, -0.5561917, -2.7552543, 0.9146824, 1.9607857, 0.4092218, -2.7102091, 1.1245851, -2.9120191, -1.9985581, -2.1078728, 1.6953103, 1.7315871, -0.2001245, 0.5898933, 0.7836690, -1.5812303, -1.1736961, 0.3256399, -0.9524814, -0.8407208, 1.0575129, 0.2472264, -2.4717003, 0.2055202, 2.8025999, 1.4438855, -2.3269164, 2.7390444, -2.5744484, -0.4991450, -2.0680159, -1.3231447, -1.9670553, 2.9790389, 2.4508656, -0.8686599, 2.3765113, 0.3431365, -0.6643942, -1.7928611, 2.4216570, -2.7884069, -1.5765209, -1.7961934, 1.3452433, 2.9110265, 1.2303118, -1.8219220, -1.4387916, 2.5074147, -1.8456955, -1.1276639, 0.5383030, -1.2412608, 2.8212675, 0.9145402, -1.3946210, 1.6005977, 2.5554362, 0.2873283, 2.7621782, 2.2780667, -0.4040796, 0.4464495, -1.8779498, 2.6803656, 1.0919362, -1.9704743, -2.9019447, -2.6692183, 2.0171652, 0.8751538, -2.4762179, 0.7833949, 0.0665479, 2.3344818, 0.8098660, -1.2708539, -0.6261810, -2.6907535, -1.7857764, -1.0337748, 2.4601973, -0.9225787, -2.3025381, -1.8113502, -2.7546028, 2.1737721, 2.3185275, 1.7100434, 1.5853766, -2.4826343, -2.0910489, 1.5161898, -0.8988345, -0.0489927, -0.4221138, 1.5278806, 0.4601884, 1.2462871, -1.6825982, 0.2356269, -1.6123932, 0.8550988, -0.2754336, -2.9683444, -2.4170893, 0.1308341, -2.2708153, -2.5513710, 1.1202680, -2.7403259, -1.4519219, 1.7862241, -1.9534082, 1.9119130, 0.7048950, 0.0738672, -0.6770710, -2.7861286, -0.1945304, 0.5879332, -2.9479530, 2.1437791, 2.6509300, -1.1527777, -2.1041240, -1.6374620, 0.4075028, -1.7220759, 1.9563895, 1.2752186, 0.1898496, -1.9707593, 0.8301975, 1.9393471, 0.5346125, -2.4889759, -2.4403356, 2.5963891, 1.4043434, 2.4241962, 2.1539612, -2.9704081, 0.3451641, 0.6184111, -2.3331418, 2.4573061, 0.9788388, -0.9684166, 1.4180670, 0.3817504, 0.7814008, -0.2887256, -0.8063817, 0.7732185, 0.7583652, 1.5345761, -2.9369207, -2.0666746, 1.1773538, 0.6854221, 2.0179621, -1.3586062, 0.0771837, -2.6375356, -1.2226113, -2.7925623, 0.1591903, 0.0698346, 0.3901696, 2.4388498, -1.3403105, -0.2446021, 2.1768460, -1.3035630, 2.3191442, -0.2795160, -1.8857661, 0.0991228, -1.1299310, -0.3068622, 1.8183242, -0.6753500, -0.5614020, 0.7393398, 2.0577454, -1.9106979, 0.4683432, -1.4348316, 0.1924204, -2.9750557, -0.2655379, 0.1693499, 2.5294182, -2.4782899, 1.1159433, -0.1615633, 1.5921848, -1.6544631, 2.4148623, 1.7454856, 0.7848833, 0.9395800, -1.8347803, -1.7452730, -1.9629272, 0.4523215, -1.0896049, -1.0953685, -1.9009616, 1.0182621, 0.4634719, 2.0026682, -1.5633717, 0.6117124, -1.3394842, 2.6810344, -2.8703054, -1.4635839, -2.8812964, 0.2163818, 1.8269235, 2.0081495, -2.6112917, -1.8021685, -2.3972419, 1.7109003, 2.6754874, 1.3119251, -1.4149269, -2.1195866, -2.5968962, -0.0408673, 0.5257302, 1.9380130, 2.5714780, -0.1910517, 2.7744617, 2.6499519, 1.6220238, -1.2991836, 0.1053020, 0.3069723, -1.3312475, 0.9751879, -2.2496038, 2.9548501, -1.8582439, 2.2766283, 1.9760078, 0.2262444, 2.0575771, 0.9251889, -0.1332939, 1.6043834, 2.6220353, -2.9797445, 2.9115192, 0.9613678, -2.8002927, -1.4581469, -1.0377567, 2.3137326, -2.3905614, 0.2651215, -2.8238030, 1.9538438, -0.8218226, -0.2868037, 1.7458996, 0.4465675, -2.7640988, -0.9651661, -1.1018883, -0.0352776, -0.4565477, -0.9355126, 2.8479599, 2.8376831, -2.4108605, -1.0590669, 2.0839101, -0.7606677, 2.9113058, -1.1215017, 0.1494032, -2.2663949, -1.2008988, 2.5577742, 2.4470562, -1.8683302, 2.8339631, 1.0940692, 0.1411565, 2.9730847, 1.0715691, 2.4969502, -0.2012309, 2.3233316, -1.4358907, 1.0153123, 0.8766342, 1.8755331, 0.4302910, -0.6877298, -0.1769293, -0.0700278, 2.4738958, -0.8846414, 1.7318973, -2.6657149, -1.0798685, -0.2116608, 0.8482216, 0.1531984, 1.7957572, -1.0834494, 0.9055639, -0.7807007, 0.4986040, 2.9761233, -2.4014165, 0.8108793, -2.6680570, 2.0672492, 0.4896273, -2.9410238, -2.6497754, 2.1570515, 0.7138747, -2.1997454, 0.0329523, 2.6184657, 0.6931318, 0.1961866, -0.2881807, 1.8025998, -1.7046810, 0.2031053, 1.2035782, 1.4471487, 0.8432122, 2.6915485, 2.8247986, -1.1444585, -1.9313899, 0.9608381, 2.3568034, -0.2887440, 0.0762962, -2.8119384, 0.9328479, 2.5258248, -0.3266954, 2.9166602, -1.5078072, 0.6026935, 0.6333275, 0.3455786, -1.1355093, -2.5627314, -0.3183445, 2.8771181, 0.7842776, 0.6820537, -1.8914184, 1.8034691, 1.6080186, 2.0685914, 0.9783015, 0.9421613, -2.2013445, -0.9547735, 0.9660231, 0.3995335, 2.0518873, 2.3041835, 2.8656644, -0.6042324, 2.8773077, -1.3175493, -0.8887908, 2.6292455, -0.7543440, 2.7924603, -0.8400863, 1.3210038, -1.7149488, -1.1151272, -2.3511033, 0.7439792, -2.2392760, 1.2774042, -0.5119403, 1.1891865, -2.5393200, 2.1352753, -2.5011709, 2.3630841, -1.6124232, 0.1646190, -2.2009859, -0.8137375, -0.5156198, 0.1943706, 1.0357535, 0.1296284, 2.9854862, -0.8675978, -1.8984936, 0.1576181, -2.4026993, -0.0829262, -1.1816254, -1.1669453, 0.8413987, 0.2489728, -1.5479498, -1.1341492, -0.2417992, 1.3035843, -0.1622541, 1.2621607, -2.0253149, -2.2939260, 2.9123313, -1.1211956, 1.9025246, 1.3323016, 2.6188349, -1.3410136, -0.0792152, -2.5649684, -2.1886231, -2.9738071, 2.6056956, -0.8215954, 1.7623715, -1.8521147, -2.3016526, -2.8235470, -2.9894598, -1.1581781, 2.4894084, 1.4694185, -2.1168502, -2.4410089, 1.9113414, 2.2349895, 1.7881586, -1.4623896, 2.5697110, 2.1764659, -1.3000729, -2.6214071, -2.5317934, 1.2858759, 1.7014427, -0.5230683, -0.5236624, -2.0597846, -1.7571240, 0.1252822, -0.8368825, -1.6104323, -2.3659168, -2.9558490, 0.8956497, 1.2186744, -1.4405914, -1.0845072, -1.4270536, -1.7629227, 1.0249317, -1.0389300, 0.9790227, -2.5412295, 0.9398306, -0.3267357, -1.8821108, -1.7236817, -0.4994807, 2.1902888, 0.4416097, 2.7047185, 0.7734643, -1.1698480, 2.4323664, 1.2967390, 2.9970495, 1.9911977, 1.0778187, 0.4825392, -0.1347564, -2.1879091, 0.9677918, 1.1192675, 2.0012550, -2.5472953, -0.0342999, 2.9918552, 1.8432018, -2.1814878, -1.3981490, -1.8549107, -2.9836133, 2.7507272, -2.5920098, 0.9293967, -0.9182083, 0.1455493, -1.0937590, -2.3801545, 1.3734389, 0.2346232, 2.9141132, 0.9092654, 1.7808393, -0.5614326, 2.8835471, 2.7166558, 0.6698291, 2.4469473, 1.1461426, -1.9722256, 1.7914399, -1.5325394, 1.1928047, 1.2622574, 2.8109631, 0.0145788, 2.1619350, -2.9039390, 2.0209792, 2.1441309, -0.3490798, 0.6683458, 1.6377594, -2.9390618, -0.1449393, -0.6676443, 0.4513642, -1.4218596, -0.0423427, -1.1580981, -1.8868823, -1.7947805, -2.5141084, -1.9105141, -0.3879839, -1.3897327, 2.1489186, -0.7781640, 1.4943134, -1.2092386, 0.4332199, 0.8065383, 2.2487376, 0.9091698, 2.2618136, 0.6885842, 2.4853959, 1.7210603, -0.2765786, 2.3321127, 2.9632710, 2.5599030, -1.7411507, 0.8364537, 2.9429951, 0.6574716, 2.9694192, -2.9854565, 1.6900069, -0.8246215, -0.3652659, -1.6420233, -1.5980035, 2.7821475, -0.0342152, 1.7023591, -0.3814957, 2.1210324, 1.5137255, -2.4665517, -0.8120593, 2.0155422, -2.4310829, 1.0920931, 2.5173831, 1.8290981, -1.8060956, -0.8577247, -1.7931687, -2.8451927, -2.6735080, -0.8611886, -1.4645985, -1.0129314, -2.7555362, 2.8125224, -1.7032590, -2.3731846, 2.5144616, 0.3252231, 0.9853244, 0.4330772, 2.3657985, -1.1487269, 1.1908465, -0.7901972, 2.5932642, 0.9765925, -1.8271584, 1.0885553, -1.4650591, -0.2132682, -2.8193983, -0.8088920, 2.9937693, -0.2979843, 1.9312420, 2.2221454, 0.4398415, 2.2159506, 2.7676346, -0.3742015, -0.7509232, -1.8096040, -1.4238979, -2.0454188, -2.3743324, 2.9927374, -2.2805380, -2.1557837, -0.5511425, -0.2644402, -1.3760140, -0.6298315, -0.3240626, 1.5880812, 0.5312325, 2.4100105, 1.3913695, -1.4322663, 0.1319617, 0.1546742, 1.0538641, -2.0603273, 2.9290994, 0.5370725, 2.5123263, 0.8733045, -1.1719780, -1.1412994, -1.9802898, -2.3670053, -0.5998347, -2.2984423, 2.4145577, 2.6722010, -0.0510579, -0.9635996, 0.4052853, -0.8366159, -0.6502491, 0.7971065, 1.7645628, -1.6442888, 2.8716308, -2.2200431, -0.1254525, -2.0067605, -2.2790566, 1.5568605, -1.0153742, -0.2599882, 2.5447521, -0.2317907, 2.1579159, 0.7499618, 1.1378918, 1.4137242, -1.6593809, 1.8493513, 0.9941138, 2.7696724, 0.8456866, -2.5494238, 1.0651606, -0.2999248, -0.3920406, 0.4353531, -0.5900873, 2.8336891, 1.8384284, 0.3686068, -2.0933811, -0.3037825, -1.4315589, 0.0027377, -1.1456297, 0.2539411, -2.5548812, -2.4022123, -1.0862711, 0.3267026, 0.9201232, 1.9721334, -0.1553948, -2.9177747, 2.4290068, 1.6525677, 0.0445467, -2.8086969, -2.9679720, -1.1525836, 1.7010071, 2.8452043, -2.6024762, 0.5900230, 2.8750062, -0.3813530, 2.3934733, -1.0643313, 2.5623713, -0.1507515, 1.8347839, 1.3363362, -2.7160640, -0.2206794, 1.5962242, -2.0134092, -1.7152933, -1.2933603, -0.4086606, 0.2588417, 1.6137543, 0.5772924, 1.3907354, 1.6867845, -1.8427954, -2.9860838, -1.0627792, -2.0700146, -0.7394871, 1.8355280, 0.3501230, -2.4308673, 1.6118396, -2.9408455, 2.3075369, -1.0527325, -1.1423548, 2.2628060, 1.0603401, -0.3865221, -1.6834122, 1.9141225, 0.2733902, 2.1709382, -0.7301674, -2.3386190, -2.9487921, 0.8003444, -1.6170643, 0.6618630, 2.1620730, -2.4660588, -1.4759390, -0.8572838, -0.5652784, -2.7120261, 0.1117577, 0.3150929, -1.3218963, 2.6064241, -1.3638313, -2.0012182, 1.2855004, -1.9863095, 1.2335874, -0.1506767, -0.5252080, -1.8419971, -0.4459362, -2.0082191, -0.4765681, -0.2209448, 1.4477909, -2.8921296, 2.8582092, -0.4093944, -2.1776744, 2.0842755, 0.5487299, 2.2134687, 1.8800279, -1.5025154, 0.4464905, -0.3145238, 2.8178712, 2.2406808, -1.5337151, -0.2781841, 1.7811769, 0.2417965, 2.5342163, 0.3305962, 1.4627645, 2.4277307, 2.3156096, -1.9637501, 2.1984628, 2.5159403, 2.6961289, 2.8098171, 1.2411738, 1.1036389, 2.1704385, -0.2085869, -0.4365357, -1.6648302, -1.0761919, -0.3796962, -1.0607764, 2.7629350, -1.8243494, 0.6787053, -0.5765959, 2.9447059, -0.1628478, -2.1529317, -0.3414518, 2.2071825, 2.2882430, 0.9916415, -1.6344449, 2.5795551, 1.9319351, 1.4091440, 1.2142884, -1.0524355, -2.8523156, 1.9071497, -2.8496023, -0.5400351, -0.1545588, 2.6211504, -0.8289387, 0.2995601, 2.9547916, -0.6074503, 1.4570902, -1.2781387, 2.2809537, 1.7200018, -1.7397199, 2.8835458, 2.6882321, -1.2098360, 1.5699560, 1.2610526, -2.3805010, 2.3213115, -1.2078863, -2.8462574, 2.9361123, -2.9102068, 1.8618695, 1.8435514, 1.2643226, 0.3184529, 1.3740391, -2.9135753, 0.7218843, -0.4831945, -2.5746059, 2.9510129, 1.2045148, 1.7001507, -0.0451061, 0.8377129, 2.5176587, 0.1859657, -2.6525824, -2.9001477, 0.8057935, 2.3823229, 0.2457998, -0.4926652, 2.9373170, -1.7653017, -1.1069599, 1.2323689, -2.3351380, 0.7817749, 1.8588568, -2.3792742, 2.1334869, -0.1156927, -1.2501091, 1.5353754, -0.5334567, -0.8711311, -0.7005431, 2.0780784, -2.0575796, -0.2802091, 1.9495938, 1.8360576, 0.6122562, -0.2716146, 1.5756510, 1.7985441, -2.9848593, 2.2619782, 0.8674309, -2.0793125, -2.0939202, 1.8247225, -2.2939749, 1.0509200, 2.2702874, -2.9955207, 0.1065131, -2.9108754, -2.3444954, 2.8336095, 2.1475924, 1.7747009, 1.4684429, 2.5600007, 2.7053124, -1.6955395, 1.5163418, 2.0626770, 0.2988213, -0.8034168, -0.5845698, 2.2128333, -0.5415805, -0.0992828, -1.9762387, 1.8182201, -1.2688550, -2.1102959, 0.8668521, -1.3393843, -0.1504119, -1.1268602, -2.6571990, 2.4152226, 1.9535645, 2.0807734, -1.8844243, -2.6750616, 2.3844301, 0.9122354, -1.8509972, 1.8539762, -2.1635874, 1.7241118, -1.6230767, 1.5329436, -1.0417966, -0.7332241, -1.1628939, -0.3684008, 1.4145694, 2.3202212, -1.1793215, 1.6668483, -1.1809875, -0.8868311, -0.6960907, -1.8378953, 2.0786010, -0.7111700, 2.4583665, 1.8489446, -1.4877366, 1.9754471, 2.7472026, -1.1124030, -1.5462028, -2.9316472, -0.0612968, -0.9170870, -2.0701961, -0.9354727, 1.4752668, 1.3351650, -2.9309617, 2.5385620, 1.8530452, -1.3486228, 0.7004151, -2.7842665, -2.1051358, 2.7384664, 1.0468108, 2.3685690, 1.5357248, 0.3601635, 0.8370112, -2.8368880, -2.9488968, 0.4496174, -1.7912519, -0.8875037, -2.0790840, 2.6544275, 1.2217982, -1.9258797, -1.0662448, 2.1236769, -1.0537595, -2.9258561, -1.8500835, 0.0373194, -0.3685569, 0.9652648, 0.6579382, 0.5735754, -0.4189056, -0.2826529, -0.8577801, -1.2858118, 0.7439400, 1.0307027, -1.0751250, 2.6891694, 0.3706900, -1.4310123, 1.3812002, -1.2827101, 1.7209388, 1.8640107, 1.2428242, 0.2424318, 2.8618024, -2.1337113, 0.5897478, 2.7459242, 0.1543271, -0.4208876, -1.2591268, -1.4213015, -0.7318079, -1.3087971, 0.2567653, 0.6642149, -1.8448265, 0.7616704, -1.5478582, 0.2732292, -1.7848982, 1.7978338, -1.3726022, -0.0296844, -0.1788379, -1.9395678, 1.3159649, 1.5696157, 1.9526549, 1.3007384, 0.2590209, 2.1569392, -0.6514665, 2.6426707, 1.0462077, 1.8650926, -0.7622907, 2.5807782, -2.2206628, -0.0523756, 2.2928411, -0.0327657, 0.5053246, 0.5231879, -2.0629685, -2.5634576, -0.6796790, -1.1941249, -1.6141237, -2.7385913, 0.6523687, 2.4414512, 1.6526913, 2.3012548, -2.6707058, 1.3522747, 2.8967400, -2.0898094, 1.9776512, 0.6657699, 1.1968666, -0.5081998, 2.7165654, 2.2204730, 0.6454324, 1.7896685, 1.8251158, -0.7424545, -0.9910009, 1.7632950, -2.7577570, -0.0964676, -2.0526622, 2.0570232, -0.9021419, 0.0074110, -0.1264903, -2.7293349, 2.7577244, -0.2843284, -2.4559699, 2.6393726, 1.7962705, 0.4086845, 0.0875447, 2.8277374, -2.5223474, 2.2007265, 2.9721267, 2.5289947, -2.6685330, 1.7064421, -1.7468457, 2.5898215, -1.6578407, 1.5492965, -1.3191672, 0.4518902, 2.0599791, 0.4743751, -2.4598416, 2.9838466, -0.9556195, -1.6580629, -2.5793204, 2.4382417, 1.3026638, 2.0794299, -1.8723906, -2.0615440, -0.1972793, 2.8433573, 1.2033883, 1.1604471, -0.7176448, 0.2442625, 1.6029338, 2.1473816, -1.0852992, 0.8640729, 1.8742029, -2.8696391, -2.5218956, -2.7227196, -2.2687173, -1.8904795, 2.8204519, -1.8749726, 2.1225633, 2.1769343, 1.8313837, 0.5759637, -1.9196942, -2.4876767, -2.8744609, 1.3948313, 1.8883466, -0.9274221, 2.0444155, 1.0558125, -1.7031227, -1.2210958, -1.7200308, 0.8986582, -2.7053576, -2.5726032, -2.2341880, -1.4551195, -2.8411452, 0.0986747, 2.9125615, 2.4185597, -1.7167749, 0.5685091, 0.2901139, 0.1630216, 1.1447992, 2.0539680, -0.6173229, 0.4875646, -1.3888233, 2.3240001, 0.0774566, 2.2700725, 2.4491782, -0.6359391, -2.0834359, 0.8621308, -0.4776596, 0.4997026, -2.3957586, 0.9871973, 2.8468504, 0.5083092, 0.5743624, 0.6287498, -2.7578971, 2.9059201, 2.7142688, 0.4204968, 2.9354537, 0.5253835, -1.5098158, 0.4710226, 0.8102967, 0.2978407, -1.9987338, -1.5352497, -2.8172453, -0.9445377, -2.0810661, -0.8034435, -0.7294693, 2.8430872, 0.1822598, -2.3558751, -1.5608193, 1.1567556, 1.8461325, 1.9906852, 0.8421484, 1.9817996, -2.5019606, -2.8236152, -1.9080595, 1.7698373, 2.2927457, 0.8382139, 1.2843581, -0.8664583, -2.6774037, -1.9295366, 1.0534660, 1.0103125, -1.4925271, 1.3489909, -0.7830498, -2.1016955, -2.4813624, 0.3560989, -1.1509657, 2.2664915, -1.5118441, 0.8798577, 2.6401151, -0.7203527, -0.1109234, 2.3990208, -2.4231368, 2.5409484, -2.6577266, 0.6053758, 1.9973182, 0.0450503, 2.3101013, -2.8040807, -0.7305345, 2.6464708, -1.5828621, 2.4597652, 0.8429633, -2.5437468, 1.0456331, -1.7615888, 0.8252650, -2.7562812, -2.8878115, 2.2512627, 0.4581093, -1.5247256, 2.3478581, -0.4715502, 1.0727651, -0.9856253, 1.2656489, 2.4055542, 2.6461035, -1.8008536, 2.5272671, 1.9795743, -2.6161955, 0.0818913, 0.7484720, -1.3155364, 1.6963326, -2.9844387, 0.5865543, 2.0540623, 1.0057556, -2.6616652, 0.0113291, -1.9837260, 0.0691968, 0.4452429, 1.6838026, 1.3200594, -2.5771805, -1.1058425, 2.3282480, -1.7322418, -2.5765498, -2.3551284, -2.9576922, -1.8352937, -2.4917617, 1.9989042, -1.3654249, 0.7093155, -1.5510189, -0.4723490, 1.9756298, -1.4449084, 0.3003121, -1.5869283, -0.0630784, -0.6673463, 0.7108110, -1.7491455, -1.3418371, -2.1694291, -2.2568286, -1.8912949, -2.0583647, -1.3582750, -1.3708235, 1.4674749, -2.9828544, -2.2536204, 2.5458074, -2.8316189, -1.3080472, 2.8522440, -1.7392184, -1.3699698, -0.1055399, -2.9105621, 1.9111560, -1.2942558, -1.8820700, -2.9763270, -2.9322751, 1.0601213, 1.7761119, -1.9416186, 0.9060939, 0.2731969, -1.2948453, -0.2025954, 2.5730738, 1.2684685, -1.7654192, -0.5609599, -0.6919241, -1.3772985, 2.8097762, -2.3072225, 0.2034328, -2.9851245, 0.0830725, 1.9149370, -1.0664587, -0.3694955, 1.4663242, -0.7899075, -0.2096035, 1.1077759, -1.6544384, -0.7754656, -1.6117510, -2.8638468, 2.7508152, -1.1419965, -0.3301882, -2.7951656, -0.9653921, -0.2571375, -2.8390454, 0.5363775, -0.5369900, -2.8563546, -0.1140510, -0.7446988, -0.8567116, -1.4180377, 1.7831481, -1.5011577, 0.1763123, 1.5217573, 2.4755685, -1.6849422, -2.4929575, 2.3838878, -2.0702608, 2.9632629, -1.4690973, 0.6751585, -2.2357885, -2.8183111, 1.7538108, -1.8110433, -0.2467183, -1.7090963, 2.2551055, 2.2066005, -2.7881238, 2.1500635, -1.3863814, 0.0801325, -1.4262124, -2.0527872, 0.8743711, -0.4027651, 1.3399882, -2.4572188, 0.2605521, 0.2855127, -1.9377880, 1.3232777, 0.4154827, 0.6402257, -0.3512390, -1.1691492, 1.0432802, 0.9727395, -1.5465813, -0.3753565, 2.5922103, -1.1306358, 2.8401169, -0.2535324, -0.2281942, 0.3223843, -1.7002352, 0.8867219, 0.2601323, 0.7725256, -1.3877158, -1.7423631, 1.9475985, -2.6831151, 1.8289042, 1.2235319, 1.5672408, -0.2402268, 2.7542684, -0.3408062, 0.8168713, -2.3749041, 1.7546043, 1.0034030, -0.2282081, 2.6066871, 2.6068815, -1.4088846, -0.5555579, 2.8646579, 0.4306410, -1.1982569, -1.0751662, -1.1707498, -1.4174288, 2.9900190, -1.3657216, 2.7588588, -1.9193823, -0.8290500, -0.5099331, -2.8276328, -0.3185254, 2.2460806, 1.7531911, 0.8098460, -0.9300338, -0.1982362, 1.5427624, 0.5225971, -2.0697932, 2.8455104, -0.3387254, -2.9929100, -0.0238930, -2.3983036, -0.1917673, -0.9698322, 1.9680605, -0.8103313, -0.9718779, -0.0533425, 1.0341472, -0.9219031, 1.2040052, -0.3732750, 1.3085923, -1.7259564, 0.8573237, 2.2652406, -0.6602044, -0.1842751, -1.8600410, -1.3132676, 2.3656129, -2.1997031, -0.3669999, 0.0767567, -1.9610973, -1.2958982, -2.4153891, -0.1528339, 0.4119860, -2.7865283, 0.0202404, -2.6067977, 2.3999056, -1.4732753, -2.4581064, 1.9679438, 1.0999643, 2.7700854, -0.8345077, 2.2546287, 2.6115473, 2.6833716, 1.6813415, -1.2120979, -0.1144573, -2.2231169, 0.8933525, 2.0059099, 0.7560344, -1.9122398, 2.6884355, -1.2396685, -1.5211786, -0.8429173, -0.7320036, -2.5125109, -1.2982640, -0.4763906, -0.8294467, -2.0616425, 2.8609734, -2.7440812, -1.2342548, -0.6083545, -1.2917791, -2.8074039, -0.2227613, 1.9298448, 1.6293656, -2.3734410, 0.6469841, -0.8263215, 0.0454834, 2.9265210, 2.0424599, 2.1827831, 0.2869029, 1.8503790, 0.5036666, 1.3492052, 0.8616955, 2.9246598, -1.8052827, 1.0588961, -1.6989427, 2.5783211, -2.9407091, 2.0293566, 2.3149326, -0.6841160, 0.4062279, -0.3714403, 0.2103661, 0.7516454, -1.0956339, 2.1469967, 1.2259600, -0.5485050, -0.7945591, 0.9961395, 0.7126064, 2.6620875, 2.9383186, 2.3074950, -2.8004412, -0.7160732, 0.1312614, -0.5031956, -1.2203061, -1.7610892, -0.5327710, 2.3364675, 0.3701399, -2.9291997, -2.7794143, 2.5265271, 0.6645864, -1.6067600, -1.2747577, -2.7283701, 0.8192705, 2.3176286, -1.5764689, -2.3866123, 1.3850920, 0.8458329, 2.2523597, 2.5866730, 1.3229146, 2.3324300, -2.9330968, -0.1994228, 1.2954288, -0.6929262, -1.2276300, 2.3369293, -2.2438678, 1.5468074, -0.7411081, 0.4973605, -2.0876521, -2.6831169, 1.3428803, -0.5151497, 0.5044558, -2.4286232, -2.3083062, -2.2685407, -2.8909092, -2.4972420, 1.7704348, 1.4783432, -1.8382060, -1.3087555, -2.9138649, -0.2312526, 2.4399225, 0.8592086, 1.2414530, -0.9609708, 0.9032829, -1.7319692, 1.3661381, -1.9818722, 0.3746582, -1.3238095, -2.2229168, 1.5366736, -0.6334204, -2.1218270, -1.9962620, -0.8256634, 2.6650610, 1.2782937, 0.8250639, 0.7501692, 1.6855966, -1.1161949, 2.0152074, 1.1989644, 0.2712566, 1.5672281, -0.7420808, 1.6976669, 0.5705824, -1.7027207, -2.7981187, -2.1092291, 2.6959571, -2.6377561, -2.7435590, 1.7654782, -2.9700596, 0.0288532, 0.8100939, 1.3573586, 0.9025364, 1.7356945, 0.3788298, 2.5328413, -1.4914978, -0.8559672, 1.9324341, -2.5750007, -0.3518815, -2.4459633, -0.5696517, -0.7906418, 2.0168149, -0.5373096, 1.1418680, -1.5044932, -0.9858097, 0.0150331, 0.9357649, 2.1757511, -2.5519519, 1.8412980, -2.2875522, -2.8511747, -2.0951767, -0.5031567, 2.8997607, -0.2131372, 2.8817370, -0.4482260, 0.2594648, 2.7892049, -0.0552679, 2.5677651, 1.9367439, 0.8169584, -1.0144586, -1.1012697, -0.6806672, -2.6300094, 0.2563362, -2.6296143, -2.9070605, 0.6883681, 1.0401348, -0.4581235, -1.8914705, -1.4181744, 2.4959750, -0.6913708, -1.2857549, -1.0331282, -2.1392737, 1.3252734, 0.5652792, -1.9127222, -1.4712288, -2.1314416, -2.9259027, -1.7752617, 1.7240966, -0.0558001, 2.1137879, 1.1895489, 2.1057124, -1.7679176, 1.3024471, -2.9187587, -2.0082592, -1.7092980, -2.7129959, 2.0727302, 0.2460285, 1.8986244, -2.7972943, 2.2268416, 2.2545789, 0.1704035, 1.1552779, -1.1856297, -0.6089014, 2.2234210, 1.8248596, -0.2664708, -2.7269643, 0.6971130, 1.2859212, 0.2944860, -2.3287374, -0.4668136, -1.2149118, -0.6268023, 1.3234899, 2.1187113, -0.0870526, -0.2551083, 2.6843244, -0.4067936, -2.7096961, -2.1631519, -2.1615341, -1.9249951, 2.2127604, 0.2643999, 2.1522655, 1.4140618, 0.1147457, 1.8581296, 1.3901385, 0.4572639, 2.0419548, 0.5768534, 2.7583303, -0.8413668, -2.6364820, -2.0314594, -1.4830227, -1.0989409, 2.8211046, -1.3781386, 0.4700680, -2.0036759, -2.7931103, -1.9440624, -2.3811585, -1.8018390, -0.5580924, 1.9842926, 1.3063329, 2.1438426, 1.4638795, -0.2886646, -2.3065319, 0.6332086, -0.5604251, -0.5307534, -0.9103982, -1.6136924, 1.3288295, 1.1844405, -0.5145992, -1.6875446, -2.2032942, 2.3349076, -2.2444827, -1.4349593, -0.8695541, -2.7292272, 0.9572045, -1.8050061, 2.8910419, 2.8442456, 0.9867765, 0.9336278, -2.1498693, 0.2741437, 2.4933028, 2.4114571, 1.8510831, -2.2558423, 1.1978109, -2.9334982, 2.9950893, -1.4360650, 0.5928946, -1.6092756, 1.5396229, -0.2349135, -1.9916375, -1.8068008, -1.8469767, -2.2188997, 2.1479047, 2.8038860, 2.2646871, 1.7725454, 0.1845193, 2.5028829, -2.0636945, 0.8079121, -0.4922575, 0.0663735, -2.7736211, 1.6917888, -0.1331106, 1.2072020, -1.7048516, -2.6959423, 0.8842196, 0.5162969, 0.5343340, 0.6603279, 0.4114421, 2.0942923, 1.8463655, 1.1526712, 0.1598658, 0.0266885, 2.5707428, -2.9126288, -2.3549700, 0.1452297, 2.3492774, 0.5199885, 2.6196456, 0.2397361, 2.1799505, -0.1568685, -1.6701414, -0.0209567, 0.4444474, -0.2846836, -1.8380434, 0.3676134, -2.4491213, -2.4082682, 1.7659272, -0.7447657, 2.6421609, 1.6454789, -2.0244421, 0.3049088, -1.7414472, 2.8123946, -2.5270487, 0.5854484, 0.8378214, 0.0449806, -0.1333212, 1.3211326, 2.0481375, -0.5923206, 2.7983877, 1.3123619, -1.6055566, -2.8046061, -1.4167368, 2.5180587, -1.2372396, -1.9086766, -0.9924344, -1.5520268, 0.9399407, 0.3794811, -0.9893087, -0.5896632, -1.5759888, -2.0034325, 0.0697662, 0.9698784, 0.0304290, 1.1914814, -1.7148604, -1.9639131, -0.2154004, -1.6426131, 0.4726983, 0.5509034, 0.1326487, -2.4756683, 2.8409180, 0.4849541, 1.0656960, 2.6744052, -2.9625314, 1.7438819, -1.7841761, -1.4770323, -1.0245589, -1.6593353, -1.9218851, -1.8889738, 0.9493583, 1.0882786, -2.6174220, -0.5981270, 0.1414073, 0.8784455, -1.4621299, 0.5314676, 2.2672452, 1.2703902, 0.1376410, 2.2445865, 1.0036056, 1.6366518, 1.4909111, -2.9593510, 2.8188767, -0.1172120, -2.2784516, 2.5578116, -1.8170748, -2.7788152, -1.2984621, 1.2323181, -1.1235460, -0.2738208, -1.2577375, 2.4498149, -1.0511503, 2.4688278, -1.1976875, -1.4074741, -2.1291158, 0.4697325, 1.9381396, 2.2311927, -0.5697472, -1.7739073, -1.4725406, -2.9521409, 1.9002849, 2.2706424, 2.3305187, 2.8941930, 0.6995840, -1.6830144, 0.9088780, -1.0937172, -1.6756112, -2.6892298, -1.4904026, 2.8072779, -2.3806429, -1.1469453, 0.5330714, -1.0197509, -0.9728791, -1.6842226, 2.6775658, 2.5475553, 1.3137924, 0.5018644, 2.5879061, 2.5410675, -2.0126178, -0.5094277, 0.3051321, 1.6205581, -0.7900410, 2.1300031, 0.3569213, -0.7711950, 0.3381163, -2.4033646, 2.4113933, -1.7493393, -2.4200764, -1.6713928, 0.9647342, 2.5144978, 2.4944596, -0.7228152, 1.6523942, -2.7332189, 2.4911265, -2.8223593, -2.4885729, 0.7389571, -0.9553738, -2.4859746, -1.6203235, 0.2954394, -0.9200482, 2.7787702, 0.2628356, -2.4263443, -1.8002772, 2.4230686, 2.1407406, -0.8033183, 2.6104895, 2.7612053, -2.5377937, -2.3169573, 1.8780457, 2.7496320, 1.8684720, 2.4010264, 0.7371540, 1.4610467, -1.5571960, -0.9373258, -0.9155709, 0.6290280, -2.8397675, -0.8896339, 0.3016679, 1.0929849, -2.1616241, 2.4000337, 2.2185850, 2.0647030, 1.9628773, 2.6143116, 1.6423320, -2.3477455, -0.7285701, -1.8069123, -2.8501723, 0.2326649, 1.7655998, -0.4387961, -1.0139296, -2.1049371, -1.6965947, -1.0949386, 2.6966676, 2.8058518, -1.8278317, 0.9671542, 0.2779216, -2.3574601, -2.6989529, 0.1889792, 0.9271327, 2.0883177, 0.5510785, 0.5393348, 2.5490100, -1.3594165, -0.0472813, -2.4574732, 1.6257403, -1.2481239, 0.8077459, -2.8584443, 2.1192402, 1.3210008, 1.8543322, -0.2111543, 2.8236513, 1.2563674, -1.4321134, 1.5344579, -0.8323285, -2.6817829, -0.2135371, 2.5892583, 0.7824692, 2.7209886, -2.8092615, 0.6045551, 2.0130957, 0.8479154, 2.1661499, -1.3277344, -2.5750351, -1.6414655, -2.9245901, 2.5844155, -2.9463202, -0.1487054, -2.5108769, 2.3433466, -2.4840291, -1.3018372, 0.7579021, 0.7870420, -1.0294452, 1.1615584, 2.5653160, -1.9628339, 1.6857889, -0.7224216, 0.5269226, -1.8382204, -2.2881081, -0.8772192, -0.8019351, -1.2270135, -0.5369647, -0.3017303, 1.1881862, 2.3969628, 0.2161541, 2.1191939, -1.5760610, 1.0454314, -0.2776711, 0.0116113, 1.3775538, 1.3265451, 1.8947193, -2.4296878, 0.7255221, 1.5782055, -0.4147288, -0.5698531, -1.1575151, 0.2235632, -0.6006033, -0.3164384, 0.6632461, -1.0780481, -1.6891931, 2.6962720, 1.1022659, -2.5844860, -2.9347675, -2.9620444, 2.5550105, -1.2252018, 0.0698074, -1.3487586, 1.1560124, 1.0016368, -1.3522835, 1.6676917, -1.1071437, -2.6599284, -1.5797484, 1.6712126, -1.2534832, 1.3495065, -0.1996030, 1.3808283, 0.8006275, -1.3801943, -1.5305734, 2.4349008, -1.1389430, -0.1511735, -1.5060133, 1.4668433, 1.3445969, -1.2721404, -0.9334931, -0.9454787, 1.9718825, 2.5310438, -0.2209738, 2.4910818, -0.6834764, -1.8053906, 2.6036291, 1.3574917, -1.7210154, 0.5750749, 1.8507795, -1.9467274, -0.2260927, -0.7294699, -2.1572496, 0.2283160, -2.0859829, 1.0685224, -2.1489844, -0.1401904, -2.4777637, 0.5433700, 1.6136671, -0.9172426, -2.8972954, -0.9519048, 1.2957665, 0.8964392, -2.8256787, -0.6380224, -2.5286782, 1.4980884, -0.9724715, 1.1786827, 1.8434202, 0.5508760, -1.9193103, 1.0309363, 1.2002173, 2.0174272, -0.6660748, 2.9386941, 0.2986273, 1.5188924, -1.1889670, -2.6984551, -2.7675065, -2.7765745, 1.1010830, 0.9917998, 2.1702986, -0.0150298, 1.5791577, 0.2747920, -1.2334004, -2.8240532, 2.0002918, 0.4045464, 0.4686324, -2.6802929, -0.2904376, -1.6553168, -2.5127216, 1.2063893, 0.1560796, -2.2345156, -1.4509625, 1.9031795, -0.3397303, 0.9319112, -0.4973973, -2.0823053, 2.6694158, 2.9461263, 0.7604430, 2.6461448, -1.3529321, -0.2094992, -1.8064986, 0.5572753, -1.8884158, -0.3634792, -2.4618812, -0.9286261, 1.4582365, -2.8454679, 0.0432023, -0.7262620, -0.5070173, 0.6565020, 1.2248492, 2.6749935, -1.1585930, 0.2569088, 2.9174619, -0.6958252, 1.1171360, 1.7655325, -1.0498500, 0.4340596, -2.2304573, 1.5128060, 1.2068847, 0.2427253, -0.0710794, 2.9022673, -2.2489619, 2.5759750, 0.2918337, -2.5914885, -2.7153252, -2.2757814, -1.3557357, -1.8004921, 1.1787679, -1.1574180, 0.3210389, -1.4966472, 1.5686408, 1.7437121, 1.1481470, -2.8908897, -0.5292702, 1.0059316, 0.2001526, 2.0824648, -2.6474451, -2.5920219, 2.8441420, 1.0215482, -1.9587196, 0.7551431, 2.6109798, -0.8884130, 0.2632468, -1.3292965, 1.1610161, -0.3313246, 1.2101142, -1.4527977, -0.2529973, 1.3423686, 1.2382265, -1.6773134, 2.9218261, -1.2739968, 0.7698736, 0.5241469, 2.6188535, -0.2541497, 0.8824040, 2.4739090, 1.4610496, -0.2811225, -1.5611040, -1.7265102, -0.7411754, 0.6456874, 1.8402550, 1.0817877, -2.1190691, -2.0148294, -1.6640528, 0.9856354, 1.4094043, 2.0682584, 0.6876083, 0.4947973, 1.5197330, -0.3403968, 1.0306441, 2.7020978, 1.0398348, 2.0263100, 1.3456951, -2.6421046, 2.7119867, -2.3568081, 0.4149698, 0.1149805, -1.3759708, 0.9098604, -0.4206787, -0.5337175, 1.1282565, -1.0864312, -2.8668264, 2.1952243, 1.1613248, -0.0673860, -1.6787316, 0.1339646, -2.2996323, -1.6421246, -1.0499550, 0.1885887, 0.0338063, -2.6183306, -2.3534297, -2.8897815, 2.5808491, 1.5059701, 1.0875996, 2.9542803, 2.3184102, 0.8249453, -1.3651835, -1.0749039, 0.2038026, -2.9266675, 2.5720964, 2.7551021, 2.6003863, 0.9639347, -1.6409875, 2.0508328, 1.7984408, 2.4349760, -1.0400961, 2.8706203, -0.5637225, 0.4175815, 1.1692462, 2.3964619, 0.8394919, -2.3310046, -2.9792603, 1.6399403, -2.7684643, -2.3899462, -2.1609919, 1.9402731, -0.8596525, -0.0871213, -0.4460283, 2.5620617, 1.3014928, -0.4041264, 0.8594226, 0.9934249, -1.0422983, -0.3501599, 0.4329727, 0.1267808, -2.3280418, 1.9745083, -0.1986156, -1.0849585, 2.9813945, -0.3958674, -0.6748159, 1.8745471, 1.0386075, -1.9445774, -0.5832601, 1.1184917, 2.2890380, -2.1533683, 0.1564705, 2.4149787, 0.0983325, 2.6245037, -2.6947762, 1.7229306, 1.8491516, 1.5289697, 1.6526286, -0.4022704, -2.0772513, -0.0206453, 1.1862265, 0.3649387, 0.1971508, -1.4899139, -1.8226298, -2.4328747, 1.8099638, 2.0868913, -1.8724177, 0.6683677, 1.7944956, -0.2416312, 1.0720109, 0.2650546, 0.8801714, 2.6947999, -1.0590103, -0.7631853, -1.8971258, 2.8563155, -0.9140186, -1.4747089, 2.0766246, 1.1387556, 1.7964485, 2.9449569, 2.8854087, 1.5561289, 1.9318747, 2.6837770, -2.2996813, -0.5312704, -0.1689105, -0.4749351, -0.4266658, 0.1489790, -1.3824903, 0.3914400, -1.2563300, 1.2821717, 0.0911681, 0.0024519, -1.3694703, -2.1822787, 2.9671916, 1.6782109, 1.6651810, 1.7953620, 2.8932230, 1.2592115, -0.0004099, 2.9800282, 0.0758289, 2.4817026, -0.7413742, 0.7370477, -2.2645835, -0.2284998, 0.1034915, -1.9447101, 2.2694557, -1.9983898, -2.7590036, 2.2735993, -1.2896299, -2.1751531, 0.0624027, -2.6571131, -1.4667214, -1.2794037, -2.7919841, 0.0359419, -0.4148895, -0.5654120, -1.0055158, 2.8775419, -1.0804933, -0.8823709, -0.8865651, -2.4188516, 2.2721720, -2.7205187, 0.1987456, -1.5411904, -0.8675275, 0.3859275, 0.8837024, -2.8566441, 1.9477224, 1.2773929, -0.1026663, -1.3969670, 2.3694790, 1.6781007, -1.0248394, 0.9196555, 2.4018430, 1.0546912, -2.3702865, -2.7062774, -2.8288986, 2.4944729, -0.4004882, -1.6590062, -2.3535963, -0.7469371, 0.6318971, 0.3371403, 2.8369300, 1.0724152, 1.5415542, -0.3281125, 1.1840022, 2.8696324, 1.0387477, 1.6442520, -1.1972109, 2.5376578, -2.6040134, 0.0050654, 1.1526993, -0.6420283, -0.4710167, 0.1789981, 1.0749018, 2.6443455, -1.1796332, -0.8892264, -1.6527535, 1.3558426, 0.6622788, -0.3677900, -1.5151313, -1.7055395, 1.6329385, 2.3582722, -0.7391464, -1.0812869, -2.9582317, 0.3321274, -0.1725444, -0.5005684, -1.7748668, -2.3630024, -1.8734890, 2.3912834, -1.2905697, -0.6729514, 0.9739264, 2.1539283, 0.1018094, -1.2918007, -2.4841996, 2.3589519, -0.8463765, -2.6855572, 2.2644104, -0.3226936, 0.0279414, -1.8879092, 2.1783359, -1.2221027, 2.9806991, -0.6665582, 2.5865782, -1.4789131, 1.7476575, -2.3239691, 1.5568208, 2.9336529, -0.9182318, 1.1130670, -0.3407502, -0.8015319, -1.9409798, -0.8731686, 1.7969460, 2.1539609, 2.2759949, -0.2256676, 1.6628799, 1.8857032, -0.2580001, 0.4168241, 2.4643207, -1.8538727, -2.9510787, 0.6500904, -1.3892282, 2.2566901, 0.5632016, -0.3292958, -2.5706287, -1.4048064, -1.3596519, 2.8484814, -1.2843858, 0.0539738, 0.3875500, 2.9124429, -2.3951132, 1.2380461, 0.8061513, 1.8216775, 1.9107133, -1.7463695, -0.8795966, 0.1719723, -0.9462170, -1.1402493, -2.4647015, -0.9368631, -2.4108788, 0.1889588, -0.2683148, -2.4292101, 1.9659911, 2.6909361, 0.9474890, 2.9162115, -1.6196272, 0.2538504, 0.0209487, -2.7257941, 2.4893946, -0.6419505, 2.0295711, -0.5084903, -1.7262967, -1.1190140, 1.5325477, -1.6563104, 1.8947950, 2.5354604, -2.3762814, 1.3575599, 1.4360569, -0.2915865, 2.6054132, 1.8921044, -1.0502901, 1.3440467, 1.8860834, -2.0768560, 1.9943836, 0.4544689, -2.1266740, -2.3140001, 1.3751911, -2.6949832, 1.7032616, -1.6140518, 1.0093192, -0.6472130, 1.1202314, -2.3026684, 2.4415909, 2.2836928, 1.4519718, 2.4502052, -2.8183591, -1.7164019, -1.8932430, -1.1115070, -1.4288013, -1.7502287, -2.1368529, 2.3183983, 1.9553708, 2.0036822, -1.4823261, -2.1855026, 0.7543864, -2.7843276, -1.1045436, -1.1545630, 2.2799700, -1.0942676, -2.1497846, -1.5104267, -2.1534897, -0.8509929, 0.9361183, -0.2051865, 2.1037959, -2.1855860, -0.7968999, 1.9681885, -1.3922168, 1.4122170, -2.8957191, -1.6957432, 2.2582310, -1.3647903, 2.5375837, -1.0055909, 1.7978272, -1.1065244, -1.8771143, -1.3030476, -0.9806063, -2.0139744, 2.9344769, -1.7813457, -0.5762509, -0.7653352, 0.3247855, 2.2124805, 0.6652285, -1.7749785, 0.3162436, -1.2359747, 0.8802232, 0.0929572, 1.4393498, 1.4077509, -2.9062622, -2.4545421, 1.4963053, 2.1298596, 1.3520789, -2.2360899, -2.5170817, -1.7204322, -0.5324893, 0.4976962, -1.0585536, 0.4484815, -2.3816757, -2.7137383, 1.0352056, 0.3417060, 0.8324133, 2.0052804, 1.8768953, -1.8536581, 0.8259330, 1.1497003, 1.7884477, -2.9359612, -0.6951613, -1.7378582, -0.5904920, 2.2799782, 1.3936917, -2.4955564, -1.4940712, 2.7145721, -2.1140465, 0.0649951, -0.3810735, -1.2494873, 2.9424350, -1.3490906, -1.6891255, 1.8797572, 1.5321115, 2.1530154, 2.0235899, -2.0635901, 0.6735616, -1.9626741, -1.9917382, -1.7591106, 0.8994820, -1.5232602, 0.9891068, -2.0103344, -0.9610179, 2.9773325, 1.4488553, -2.3761333, 1.2647832, -2.6533800, -0.2246688, 0.6801636, 0.4741215, 2.2965509, 2.5405495, -1.9305077, -0.0171405, -0.2614862, 0.8245159, 0.1610389, 0.2518784, -1.0204004, -0.0111499, 1.5918429, 2.8102683, -0.7315727, -0.9023423, 1.7519760, -1.9167747, 2.2367203, -0.0426625, 2.4513946, 2.8742536, -1.4524389, -0.1115864, -0.0337808, 1.5641894, -2.1374891, 2.3394541, -2.4910297, -2.3736973, 0.2209650, 0.3458578, -0.5005771, 1.5614608, -0.6307671, 2.6636051, -0.1405854, 2.7316020, 1.0366162, 2.9418266, -0.1429010, -0.9675913, -2.9573177, -2.9434267, -0.3731679, 0.1067155, 1.5775927, 0.9432656, -2.0919523, 0.1662257, 1.0727488, -1.1042745, 2.7689285, -1.1635115, -0.7740340, 2.1366532, -0.5120563, 1.7932125, 2.7143831, -2.7691796, 1.0888875, 2.6523738, 2.2407927, -0.4414625, -1.2009725, -0.4106058, -0.6275878, -1.9312175, 0.8658490, -0.7058895, -2.8894322, 0.8044130, 2.6929670, -1.5168462, 1.1598375, -0.5195148, 2.6875938, 1.0087141, 0.2423690, -2.3632173, 1.6411540, 1.5978333, -2.3160699, 0.4556444, -1.9754069, -2.0110125, -2.0311330, 1.3194541, -0.0490528, -2.5803440, 1.9423533, 1.1698608, -2.1971197, -0.8266906, 2.4050886, -1.0457988, -2.8283474, -0.3619271, -2.1251539, -0.7185260, -1.1936631, 1.4587760, -1.8526359, -0.2442774, -1.0507360, 0.6643322, -0.6468434, 1.1007906, -1.3172159, 1.4958873, -0.4185608, 2.2554517, -2.2144080, -1.5183857, 0.2287259, -2.0824601, 0.6806877, 0.5239830, 1.6213139, -0.5295686, -0.6123455, -0.3299208, 2.9627587, 2.1609544, 0.7306745, -0.3536996, 0.8648042, -0.0107556, 0.5563253, -1.4150572, -0.8727354, 1.7045240, 0.2422660, -1.9675813, 2.3998704, 1.2408928, -0.8462677, 2.5386144, 0.8989565, 1.0722134, 1.4754168, -2.6578095, 0.7917410, 0.2518352, 2.7770565, -1.6927019, -0.9069547, 0.6937956, 1.8118292, 1.4657977, 1.6499550, -1.9093678, 1.6016672, 2.9462244, -1.5291002, 0.8729590, 1.6649800, 1.8471859, -0.0921219, -2.6374733, -2.7870960, 1.8837198, -2.0499895, -0.4946272, -1.0308865, -0.1609454, -0.1261321, -2.5382789, -0.3218134, 1.8543531, 2.2648123, -0.3317457, -0.7465101, -0.4652393, -2.6359527, -2.9831871, -1.8001781, 2.4441152, -0.4254941, -0.9714003, 1.3048707, 1.9364892, 0.1989429, -1.3276407, 2.5982068, 0.8736684, 0.5124597, -1.9403549, 0.4400453, -1.8829024, 1.4911714, 0.4730502, 2.4722706, 1.3535375, 1.2369254, -2.1041016, 1.1254182, -1.3134398, 1.1766882, -2.2733701, 0.8459110, 2.2576526, -0.5385826, -0.6113111, 1.9070254, 0.8045966, 1.1241913, -2.3495071, 1.7460611, 0.1448644, -0.1904890, -0.4045659, 2.7795005, 1.4751990, -0.6674187, -2.5507093, 0.2030538, -0.2692014, -2.6217253, 2.7209130, -0.0345736, -0.6282908, -0.8736098, -2.4026508, 2.1056605, -1.2177200, -1.7237630, -0.4934834, 0.1289675, 1.7176823, 2.6431999, -2.8293549, -2.6321991, 1.2287625, 1.0290202, 0.6316410, -2.8051481, -1.1754169, -0.1512916, 0.4032677, 0.5490186, -0.6788442, 1.9478857, 2.0590555, -1.7040275, -0.8266720, -0.5077819, 0.5894257, 1.4900348, 2.3215805, 1.8013488, 0.3438201, -0.8274180, -1.6088323, -0.3611190, -0.4598206, 2.9183847, 1.9363682, -2.3514224, -2.2227259, -1.6925201, -0.5801150, -0.7014093, 1.3379582, 1.3345020, -2.6102805, 1.0340657, 0.0950508, 2.7118344, 2.2549243, -1.7944578, 0.8886559, -1.6920553, 1.8236820, 2.4413825, 1.0226802, 0.8347702, 1.3612298, 2.0169374, -0.0753581, -2.5647480, 2.5113865, -1.4995078, 0.0460619, 1.8805909, -0.9555030, 1.6477782, -1.3508497, -0.5109600, 1.7161824, -1.9356188, 2.8784849, 2.1395209, 2.5442767, 1.5916446, -1.9272739, 0.4771991, -2.5477749, 2.5653464, -2.6951755, 0.7098542, 2.6758043, 0.2559537, -2.2485367, -2.6685046, 0.6916883, 1.9410004, 0.2091923, -0.4386480, -0.7369906, 1.3450719, -2.3366159, 1.8566166, 2.5931245, 2.0692529, -0.1774360, -1.0984693, -2.6529387, -1.8842363, -2.5040193, 0.8633573, -0.5938961, 2.5152711, 0.9716124, -0.6287754, -1.7735882, -0.7446117, -1.1069206, -0.5352360, 0.4325741, -1.6197771, -1.9263385, 1.1817253, 1.5157346, 0.5527270, -0.4255365, -0.0006920, -1.0274411, -1.8450064, -2.1935538, -1.3004155, -0.4128389, 1.5186578, -1.5064052, -0.3992769, -2.8860171, -0.4211497, 1.6081145, -1.0839095, -2.3088657, -2.5115435, 2.2794044, -0.3706322, 1.3227494, 0.2703471, -0.5612499, 1.5913938, 0.9805876, -2.7110857, -0.4797490, -2.8291773, 0.8045318, 2.2173060, 2.2878503, -0.2371392, 0.3249561, 0.5830039, -0.7491246, 0.7867096, -2.4699055, -1.5524765, -2.4647461, 1.7322005, -0.6696453, 1.9075731, 0.7549530, 1.7624442, -2.8692598, -0.6889116, 0.9746551, 0.2208775, -2.4180421, -0.7243910, -0.7207610, -1.5957735, -0.1000400, -2.2506119, 1.4959637, -1.2871287, -0.1025470, 0.1829531, -2.5310866, -1.0562694, 0.4305466, 1.1116550, -0.1867656, -0.9307736, -1.9929554, -0.5467123, -2.3586867, 2.5430691, 0.1858240, -2.2750922, -0.1376593, 0.6767229, 2.0055602, 1.1808723, -2.7447532, 0.8980540, 0.0772440, -2.0398544, -2.7438451, 1.6259597, -0.9553521, -0.7801304, 2.0049282, 2.9398424, -1.0702306, -2.1168996, -2.0416170, 1.3785923, -2.5926850, 1.0390946, -1.1574019, -0.7132420, 0.2734655, 1.3967249, 2.4575069, 1.4214275, -0.0668784, 1.3928680, -0.4120073, -2.7979377, 2.6651927, 2.7760301, -1.8485916, 0.1390376, 2.6033872, 2.3731228, -1.7451586, 0.8325962, 2.3761913, -1.5268622, 1.7894355, 1.2926317, 2.4120051, -2.9943664, 1.5151347, -2.5051500, -2.6444565, 0.1493495, -2.0373937, -0.0515417, 2.2976269, -1.3238267, -2.9406643, -2.7537111, -1.0604598, 0.8613906, -2.0844975, -0.0685212, 2.0613430, -0.9591255, 1.1293803, -0.7282211, 2.2175269, 2.4242548, 0.8512171, -2.3346040, -0.6742826, -2.5614914, -0.0130313, -1.6337592, -1.8547938, 1.6781894, -1.8701950, 2.6305676, 1.0458117, 1.4097527, -0.3030116, 0.1706202, -0.0997305, 2.9243656, -1.3471538, -2.7494799, 0.9894578, -1.7116989, 0.4116193, -0.8716717, -0.0325625, -0.5310757, -2.0841364, -1.8789701, 0.6990849, -1.5842051, -2.6421534, -1.9632266, 0.0472854, -2.5241316, -0.4943429, 0.1470748, -2.6732500, 2.0138913, 1.9013081, -0.7417802, 1.4396681, -2.2319511, -2.4684710, 0.9345021, -0.9673472, -2.7694178, 0.5690039, -1.5052723, -1.5785337, -1.0897557, -1.3056671, 2.9203166, -1.7758468, 2.6161321, 1.4677514, 0.8884222, 1.1094984, -0.0578506, 2.5794072, -2.8453195, -2.9410432, -1.4636468, -0.4812051, 2.0318668, -0.9069256, 0.7700721, -1.7329202, 2.7328775, -2.9528846, 2.3844544, 0.5625010, -1.2629683, 1.6787202, -1.2234445, -0.6106854, -1.8477321, -2.5704755, 0.7858727, 1.0341762, 2.5851653, -0.2452754, 2.7613799, -2.6940972, -1.2159570, -0.7063653, -1.3779938, 1.8720782, -2.5275128, -2.0654881, -1.3038211, -2.4652363, -1.1270873, -2.1256460, -2.9914899, 1.8846489, -2.4404785, -0.5126766, -2.8117912, 2.5900067, -2.5923891, 2.8501839, -1.9304444, 0.2033321, -2.2504419, 1.4925323, -2.9500139, -1.3922348, 1.6349420, 2.0449034, 1.7383640, 2.0677755, 0.2452044, -2.4821752, -1.7241185, 0.1891097, -2.5512692, -1.2766243, 2.7032303, 2.0594200, 0.5038068, 2.9359277, 0.4792132, 0.2217329, 2.0401450, 0.9586963, 1.1161192, 2.6023374, 1.9791698, -0.0160477, 0.4282678, -0.4256023, -1.4846920, 0.3257271, -1.3356290, -1.4922830, -0.5841838, 0.6646986, -0.8536927, 0.9543134, 1.1195122, -0.8371800, -0.4028238, -1.4547128, 1.2306021, -1.4179080, 1.9255175, -2.4631044, 1.7002114, 2.9943265, 1.5694730, -0.4246447, 0.6873153, 2.5256696, -0.1803972, 1.3017915, -2.8728148, -1.9913368, 0.3396982, 2.2304179, -1.9865419, -0.4319300, 2.3424087, 1.4413776, 1.6222765, 1.6235918, 0.5569569, -0.0089463, -0.0956309, -2.5100063, -1.8787572, -2.7184046, -1.9358166, 0.7386632, 2.6771919, -0.7123779, 1.1437926, 0.8210358, 1.4300204, 2.2206613, 0.7998181, -1.1064798, 0.7351197, 1.9705326, 2.4720239, 1.6906173, -2.4013767, -2.3493172, 1.8080084, 0.9508681, -2.0578745, 1.0356559, -0.1402811, -0.0951342, 2.5867359, 1.9537267, 0.0392803, 0.3871637, 0.3527258, 0.7576648, 1.4197035, -0.0151841, 0.7506823, 1.0906425, 1.1608549, -1.8603324, -0.4505152, 1.9362832, -1.5389217, 1.0650490, -0.7252602, -1.4728714, 1.8775472, -0.2296435, -0.3072488, 1.1724754, -1.6757912, -2.3079057, 1.0504699, -2.0819913, -0.9674736, 1.7811321, 2.4198991, 1.9606676, 1.7131432, 2.4777274, 1.1861515, 0.3224512, 2.6746817, -1.1585997, -2.4805994, 0.3183342, -0.7560267, -0.3013422, 0.0370007, -0.1201556, -1.0747571, 1.2244132, -2.8129453, 2.4159154, 0.7767780, 1.5164903, -1.5278360, -2.6134863, -2.6279116, 2.5568834, 0.1311238, -1.3508781, -0.2330924, -0.6013837, 1.1767107, 2.3271863, 0.0970165, 1.3980686, -2.2584791, -2.6101869, -0.7449564, 0.4994273, 2.6127898, 1.0511579, 0.1972315, 1.9911316, 0.2242351, -1.2519555, 1.4642125, 2.4550977, -0.2664855, 0.6366780, -1.8333734, -0.9785470, -1.3776121, -1.2519539, -1.4613658, 2.7517760, -1.4644457, 2.6353145, -2.3399311, -1.0098588, 0.5789256, -0.0255538, 2.8470338, -0.9017638, -0.1068883, -2.6378680, 0.6243256, -2.6210253, -2.3329380, -0.9272802, 2.4540008, 0.4191707, -2.0345299, 0.7544554, 0.2131334, -2.1841153, 0.1785419, 0.4181768, -0.8432541, 0.5277870, 0.2974365, -1.3460967, 0.7204510, 2.5884003, 0.2821836, 2.3958907, 0.7231284, 0.0650873, -1.6860096, 0.6566120, -1.3402215, 0.2204201, 1.7253816, 2.9077322, -2.1117129, 0.2275158, -0.2371496, -2.3832028, 1.9442344, -1.2291940, -2.0293144, -2.8315288, 2.3858388, 2.4489611, -1.5138199, 0.1517202, -2.7135367, -1.3286428, 2.6979218, 1.2594799, -0.7910451, -1.1066100, 1.8046372, -2.8139491, -0.8969320, -1.9809114, -2.4191667, 1.1946921, 1.6507736, 0.7950459, 2.0576455, 1.8020493, 0.5389994, 1.5924049, 0.9181959, 0.0697358, -0.3594174, 1.0726308, 1.0808109, 0.6562864, 0.7561583, -1.6409176, 2.4685848, 1.2381941, 0.3960441, 1.5286791, 1.0868504, -2.0699569, 2.0799829, -0.3232925, 1.4528518, 1.7440543, -1.7781581, 0.6488502, -1.4723385, -2.6355891, -2.1567801, 0.1053335, 0.1852978, 1.5779263, 2.2734339, 2.5119967, 2.5675381, 2.1252138, 1.5136475, 0.5624561, 1.6699814, 0.7043991, -2.7956257, 1.3890359, 1.2846648, -2.9567038, 2.3157683, 1.3543212, -1.2813881, 1.3293518, -0.2054878, 0.3350399, 0.9901608, -1.7680799, -2.8931328, -0.7080173, 0.0589902, 2.0004146, 1.6022610, -1.1391519, -1.9729754, 2.1602098, 0.4287585, 2.1244229, 2.2273216, 2.9446939, 2.0101983, 2.8430189, 2.7768658, 2.4938386, -2.1529353, 1.6068259, 1.5241928, 1.2005206, 2.4702329, -2.4603307, -1.2792345, 0.1389811, 0.2947822, 1.4342956, -0.9773418, -1.2160389, 0.6666885, -0.9517086, -1.7169715, -1.4546749, -0.7354775, -2.5203226, 1.5270202, 2.6805747, 1.4467756, -0.3184058, -1.3979394, -1.7181460, 2.8663034, 2.4224627, 0.3159663, 1.1681837, 1.7505577, -1.0540509, 2.7435352, 1.1176091, -0.9438068, -2.7228308, 0.4540646, -0.6692979, -2.3128386, -2.1583480, -1.9458854, 0.6169611, 2.4761246, 2.7338699, -0.9783063, -0.2154977, 1.5536672, 0.5792992, -2.2523444, 1.4179318, -2.1651964, -2.1360809, 0.6297456, -2.7593438, -1.8385471, 0.4390709, 2.4636268, -2.0884041, 1.3402412, -1.5487623, -1.5425371, 2.4212514, -2.9943274, 2.1771449, 1.1747888, 0.6076876, 0.6557948, 1.0158448, 2.9831179, -1.5819440, -0.5242162, 2.1767828, -0.3128429, -2.9144030, -1.3114079, 2.1906147, 2.1112061, 2.2442529, -1.9983339, 0.1156998, -1.8924436, 1.5943900, -2.5990841, -1.2849910, 0.1616793, -0.8476348, 1.9128135, -1.1821586, -2.3928171, -2.1474731, -2.5316257, 1.0602172, 1.0337591, -2.9133754, 2.9269145, -0.4936134, 0.7414270, -2.9613635, -2.8390568, -1.0072504, 2.4713025, -2.0964645, -0.0454044, -0.3731113, 2.2123210, -1.1434951, 2.9163429, -2.2469878, 0.2200340, -0.8263998, 0.2289010, -1.6770205, 0.8381352, 2.8176167, 1.0498123, 2.0576354, 1.4023614, -0.1381644, -0.1252577, 1.3247484, 2.5922736, -0.2778088, 1.9959282, 1.9320127, 2.4483298, -2.8119544, -2.8411717, 1.0070857, -0.7279842, 0.5166012, -1.9092448, -0.8770331, 1.2288802, 0.8464884, -1.7913210, -1.7995877, 0.6250318, 1.6069269, -1.6330905, -1.3394804, 0.7219097, -2.8823360, -2.7134405, -2.9912427, -0.0746364, 0.6150895, -1.4942205, -1.5752316, -2.4934232, 2.6103250, -2.9869983, -1.6025418, -0.4396260, -1.6260243, -2.4966483, 0.7481000, -2.0465925, -1.9146622, 1.8339351, -0.1138441, -1.6991243, 1.6380141, -2.9643933, -0.1159944, 1.7969160, -2.9256233, -0.9882193, 0.2795916, 2.6718566, -0.6763195, 0.7237665, 0.3217816, -1.2267966, 1.4301360, 0.2543050, -2.0177207, -0.4432968, 1.1997924, 2.7155361, -1.4915216, 2.9253556, -2.9563903, 2.6567566, -2.9624302, -2.7198583, -2.7939154, -2.9753752, 2.6686465, 1.2337032, 2.3226727, -0.6032942, -2.6710755, 2.2622624, -1.7090637, -2.3882325, 1.6797622, -0.0301304, -2.0227944, 2.5327229, -1.5613255, 2.0236975, -1.0351895, 1.3502886, 0.4575648, 1.6815330, 1.5684237, 0.1107819, -0.9096126, -1.9795333, -2.7488899, -2.3859125, 1.9261755, 2.3533089, -1.5704912, -1.9260879, 0.7484132, -2.5803128, -1.7775928, -0.3527641, 1.5616242, -2.2647986, 1.5672011, 2.6305416, 2.5920888, -2.3910170, 2.1460191, -2.9813728, -1.7314653, -2.5300958, -0.6480946, 1.1395040, 2.9523720, 0.6262421, -1.4078439, -1.1475230, -0.9482321, 0.4622595, -0.8447258, 2.9223331, -1.3249990, -0.8124064, -1.8033663, -2.0145743, 1.3212688, 2.5692527, 2.7943714, 1.0720738, -1.5700753, -1.8362480, 1.0430671, -2.2832940, 1.8451702, 1.3025234, 1.1496870, 0.6185796, -0.0240178, 0.9515752, -1.9289805, 2.9877216, 0.2191507, 1.1269093, -1.8602446, 0.7527767, -2.3128837, 0.4271805, -1.5612495, -2.3409141, 2.4629432, 1.8618237, -2.1263927, 2.3395088, -0.0765445, -0.5821758, 1.4542050, 1.4069796, 0.7942523, 1.7198090, -0.8742714, -2.0515206, -2.1393170, -2.8145044, -1.1351348, -0.3610599, -2.9604500, 0.8635343, -0.9616761, -2.0176324, -0.4981394, -2.1162554, 0.5105758, 2.8691310, -2.2764248, -0.5595060, 1.1661863, -0.4900028, 0.1688583, -0.6903034, 0.9144493, 0.5237892, -1.8439340, 2.7207143, 0.9570627, 0.3382306, -0.7632022, 1.3092409, 2.9204649, 1.8582604, 2.3075137, 0.3782695, 1.9356775, -2.6129667, 0.5020823, 0.8470648, -0.2877516, 2.6285079, 1.4953637, 2.0980395, 2.6794553, 2.1306104, 0.8995583, 1.3563450, -0.0664813, -1.1265710, 0.2566990, -2.3765097, -1.4268553, -0.7278489, -1.5187537, -1.4612712, 2.8520545, 0.3487226, 2.0089191, 2.2290274, 1.6936494, -1.8538784, -0.1525317, 2.9372055, 1.5399349, -2.6755948, -0.7354602, 1.7105238, 2.8917153, 1.3430876, -0.2488672, -1.6465223, 1.1422599, 2.5891537, 2.9478575, 1.5250615, -0.3427170, -2.9007160, -1.6266121, 0.0088667, 0.0800767, 1.4107517, 1.5132156, 0.5423988, -1.0013136, -0.7373925, -0.0824629, 2.5128762, 0.4141175, 2.0636659, 1.9287245, -2.3236154, -1.5027373, -2.1796979, -0.8312790, 0.3037361, 2.1079695, -2.9168071, -1.5822629, 0.3229404, 1.8527595, -2.4633541, -0.7595892, 0.1492531, -2.9604665, 2.6274724, -2.5541728, -2.1960779, -0.6548288, 0.9323413, 1.1847380, 2.4807662, 2.2309652, -0.7180121, -1.7218763, 1.7704366, -1.5928659, -2.7414276, -1.7370882, 1.5761903, -0.5225891, -2.1271784, -0.9448735, 2.6234764, -1.2165242, -1.7494884, -2.8047693, -0.0292116, 1.0547753, -1.4575132, -1.3930879, 1.8352372, 1.4753862, -1.3835359, 0.7085792, 0.7326964, 1.1649280, 0.1098104, -0.5146073, -0.5539026, -1.9569064, -2.7192358, 2.9889935, -2.8309225, 1.9873359, 1.1594913, 1.6535363, 0.6550989, 1.2319942, 0.2754955, -1.7375855, 1.7432973, -1.6725076, -2.8417370, 0.0247126, 0.6801791, 2.4012191, -1.9731452, -0.8414916, -1.5652772, -1.9710613, -1.2263543, 2.9261207, 0.3256376, 0.4920433, 2.9528342, 0.1422812, -0.9643146, 2.9870621, -0.9874027, -1.6665130, 2.6215618, -0.8317672, 0.3609345, -0.6012590, -1.4569081, -1.0487993, 0.2255016, -2.6316194, 1.9495046, 2.1938144, 1.0478005, -1.0368773, -0.4049171, 1.0665002, 1.8470732, 1.8305455, -2.7596019, 2.6606894, 1.0800696, 2.8906324, -2.0165279, 0.8781187, 0.8741900, 1.7987329, -0.3957045, 1.7482102, -0.9367998, 2.3200296, -2.8270043, 1.0839189, -1.8452330, -0.9518633, -1.8263326, 2.0230787, -2.4806369, -2.8099271, -1.7706231, 2.8895067, -0.6726223, -1.0248627, 2.7106785, -1.0082413, 2.0894818, 2.2648872, -1.3012480, -0.7536116, -2.0789771, 0.6951624, -0.0992962, -2.2802300, -2.0413623, -1.5007342, -2.2068135, 1.3712549, 1.1260024, 0.0797329, 0.9953381, 2.1667766, 2.9000574, -0.0861247, 1.3356928, 0.9292654, -1.3605494, -0.6385973, -2.5772347, -0.6496099, -0.6822974, -0.0030114, 1.1784882, -2.4366380, -2.5236719, 0.7240618, 2.7251474, -2.5993238, 0.7892850, -2.7502414, 0.8146159, -1.1905411, 1.7165819, 1.5822982, -2.7096877, 2.5990128, -0.0145802, -0.9755537, -1.9864763, -2.7036628, 0.9945190, -0.2788020, 1.5601044, 0.9265302, -0.3084860, 2.0386146, 0.9882662, 0.8410817, -0.4694067, 2.2472006, -2.7328041, -1.6870877, 1.0512815, -2.7313614, -1.6054064, 1.1565029, 0.3482166, -1.4567974, 0.9865063, 1.0934233, -0.9808005, 1.9430768, 2.3342066, 0.7781535, 0.9788652, 1.0187933, -2.8085644, -0.5025205, -2.6636854, 0.8330482, -1.5719949, 0.4931525, 0.9627076, 1.8942991, 1.9246273, -1.3893339, -1.5850160, -2.8456102, -0.2590670, 0.0241291, 1.2145132, -1.7147631, -1.1090574, -2.2923959, 1.8376368, 1.3154051, 1.2471854, 1.9335377, -1.8634069, 2.9568108, -0.3716599, -2.0259255, -1.7317291, -1.0623009, 0.9393323, 1.6714617, -1.7635129, -2.1462233, 0.8708822, -0.5368493, -2.0561552, 1.8944607, 0.1597335, -0.2404044, -1.6333906, -1.9963300, 0.8683341, 1.0216861, 2.9771490, -0.1348256, -1.2063377, -1.1501009, 1.0790666, -1.5337711, 1.0090484, -1.2487039, -0.1127489, 0.0574801, -1.4278137, 2.3272467, 0.5837185, -2.5833496, 0.2342355, 2.1547140, 1.8870283, -2.0099986, 0.6310067, -0.9638803, -2.7837276, -1.4877928, 0.3441679, -2.5031214, -2.7207024, 1.2927608, 0.9710515, 2.2462752, 0.7233333, -2.7244101, -1.7079876, -2.2500971, 0.7399123, -0.7388021, -0.8180460, -0.1541326, 2.7187128, 0.2788272, 0.2114331, 0.8945514, 2.1896248, 1.9271862, -0.7307687, 1.9386922, 1.2322866, -1.1017456, -0.3487095, 2.5010391, 0.1911470, -0.1120439, 1.9048201, 0.9863319, 2.3157479, -1.8557647, -2.8726068, -0.7144961, -2.0277188, 2.2110567, -2.3156594, -1.3869185, 0.5647291, 2.3912793, 1.5031933, 1.8634769, -2.9395758, 0.9064631, -0.0465871, -0.8397804, 0.0151774, -0.6716056, 1.7621311, -2.3605577, -1.0053672, -0.0210941, 0.4782855, 2.8176531, -0.9404110, 0.1141604, 1.9818238, 1.0668255, -1.2280843, -1.9334220, 0.8335752, -1.5284786, 0.9286313, -1.4532219, -1.0743614, 2.2035467, -1.0244209, 0.4524791, -1.4198160, -1.8475322, -0.6007970, -2.8086697, 1.6439996, -1.4681064, -2.6377254, 0.5657356, -1.7456060, -2.1018656, 2.8168153, 1.5327052, 1.3557180, 1.4777876, 1.0251620, -0.9834132, 2.1458915, 2.5128371, 2.7137593, 1.3509308, -1.6136117, 0.1325019, 1.3441331, 1.6121391, -2.7924737, 0.4916447, -2.3137470, -2.7848982, -0.7539787, -0.7757549, 0.7977458, 2.5196707, 0.2164295, 1.4132255, -0.8239160, -2.1679258, -1.1789784, -2.7320671, 0.8172988, 1.1206406, -1.4262843, 2.1152431, -2.4526066, -1.8688534, -0.5073304, 1.3273777, -1.2861214, 0.6718110, 0.8981626, 0.5060007, 0.6785249, -0.5185401, -0.9143499, -2.4297972, -0.7427988, -1.0906686, 1.0590956, 2.5512235, -0.1521870, 0.5238273, 1.3357581, -2.9465626, -1.5641982, 2.3129222, 2.9033436, 0.7224817, -0.6641415, 0.4944516, -1.7313599, 0.1826410, -2.3793119, -0.0165791, -1.8099073, 2.9001312, -0.3801332, -1.1391284, -2.8021860, 0.9260575, 1.7532860, 2.3597246, 0.0583827, 0.9575774, 2.1946098, 1.0557186, 0.3632254, -2.7260005, -2.8667138, 1.7380930, 2.8765011, -1.0654563, 1.5951050, -0.3011768, 1.1611062, -1.5077208, -0.7250073, -1.2131459, 0.8252430, 2.0157391, 0.2732854, -2.2574970, 0.6080738, 2.9697753, -1.4866057, -1.8125294, 1.4225773, -0.8099765, -1.2790249, -2.9133621, -0.9798591, 2.5401327, -1.3994812, -2.8482290, 1.4009607, 0.6440566, -0.0881436, -2.2265096, -2.6358205, -1.8510079, 0.7577829, -2.9047972, 0.5694009, -0.1248517, -0.7485144, 2.9659904, -1.5647706, -2.4475029, 0.6205009, -0.7005075, 1.2271329, 2.2897045, 2.8402924, -2.4773290, -1.0565600, 0.7538679, -0.2968332, 0.7030878, -2.3410934, 2.2881827, 1.9963076, 2.5786977, 0.9341983, 1.3867988, 2.5376485, -0.0423620, -1.0103831, -2.8328037, -2.8958100, 2.5247765, -1.4505308, 0.4198141, 1.8244588, -2.0702264, -1.9231865, -0.1604105, -1.4758346, -2.0295263, -1.0032046, -1.5283908, 1.4389132, 0.8665983, 2.8220219, 2.9331439, 2.5789314, 2.4190159, 1.3577563, -0.1053213, -1.2426670, -2.5773538, 2.3540017, -1.1498071, 0.7753672, 0.2072255, -1.4531528, 2.8641035, -1.1971309, -2.6191845, 2.9063073, -0.0450908, 1.7277749, -0.4319434, 0.5187176, 1.2259523, 0.3790746, -1.9521823, 0.2379017, -2.5148859, 2.2773292, 2.0867761, 0.2501841, -1.9111912, -2.7021212, 0.6985916, -2.6058813, 1.4570822, 1.5059125, -2.6682442, -0.4486553, 0.5296342, -2.2083631, 2.4918160, -0.2019975, -1.4653366, 2.6714460, -0.7394957, 1.5151877, 0.9473406, 1.7446577, -1.8359983, -0.0034084, 2.9874980, 1.2525770, -0.6114602, -0.1351516, -1.8772852, 0.0333585, -2.1532100, -2.9858631, -1.9156199, -1.7762967, 0.4810657, 0.2731672, 0.8353681, -0.0239810, -0.7848465, 2.4525829, 1.5844366, 0.7775841, 0.4704033, 2.3867158, -1.1036819, 2.5401483, 2.2960970, -1.6180077, 1.8757254, 1.6948931, -2.7125149, 2.7689038, 0.7585525, -2.7372075, 1.6756445, 2.9846808, 1.6380267, -2.6500161, -2.7263904, 1.5481572, -0.7318222, 2.0983924, -2.6248315, 0.2988894, 1.1831656, 2.0417642, 2.8073981, -2.9001361, 1.9891103, -0.4872648, 1.9040536, 2.6837978, -2.0041785, 0.9850764, 2.9819866, -1.1572081, -1.5400224, -0.0171987, -1.0213449, -0.5816555, 0.7064418, 1.6238504, 0.8715284, -1.2352366, -1.0683733, -1.2476769, -2.4680943, 2.9708698, 0.2230209, -1.5653560, 0.0292373, -1.7771650, -1.9823033, -1.0220443, -1.1920262, -0.3020521, -2.5752950, 0.9653428, 2.2563952, -1.9970893, -0.5061781, -2.5182596, 2.4604912, 2.2559172, -0.1500541, -0.8061987, 1.8862678, -2.8240897, 1.0201338, -2.2660666, -1.3089319, 1.7156447, -0.1534503, -0.4594935, -0.9321401, 1.0907786, 1.7078927, 1.1942217, -1.9252083, 1.5711110, -0.1807472, 1.9737335, -0.7362138, -0.4373959, 2.3745196, 0.8188940, 2.4264595, 0.4286129, -2.5813692, 0.9198657, -2.0264455, -1.8325156, -0.2153014, 2.3699933, 1.1267198, -2.3897631, -2.2409915, -0.3459683, -2.2308153, 2.3960800, 0.2934987, 0.3852452, -0.3846697, -1.9159654, -2.0461001, -1.2260260, -2.3601156, 2.8759282, -0.9638342, -0.0636866, 2.1610389, 1.0514992, -1.7158630, -1.4566643, 1.4334064, -0.8454233, 1.9436244, 0.0705983, -1.7534019, -1.4151513, -2.3489959, -0.3489684, -1.5821723, -1.6095886, 2.0773892, -1.5448042, -2.2660495, -1.3090968, -2.9532824, 0.4497670, -0.5059318, -2.8271314, 0.0367679, -1.0489132, 0.5247005, -1.7327810, 0.2169870, 1.1690485, -1.6468392, -1.2412470, -2.9978692, -1.7492706, 1.3012010, 0.1184864, 1.5131942, -2.5881241, -0.0855265, -2.1384913, 2.7954950, 2.2794679, -0.9193915, -2.1517246, 2.2431840, -1.6935083, -1.8405548, -0.8753732, 0.5521554, -0.4166712, -1.2822242, -0.5837516, 1.0730054, -0.2433895, 1.0178278, 0.4966163, 1.3702224, -2.2520963, -2.4899451, -2.4027284, -1.6615509, -0.7060132, -1.7460305, -0.0439235, 2.5573767, 2.7884397, 1.6295932, 1.8865269, -2.5864131, -2.0500739, -0.4900841, -1.1732292, 0.3184292, 2.1157396, -2.4114227, 1.1948997, 1.1598677, 0.5738076, 2.8843175, 2.0419706, 0.1235445, 0.5814506, 2.6008974, -1.8974137, -1.7088389, -2.8783539, 0.8736214, -1.2913917, -2.4985147, 0.4018654, 1.1875748, 0.1425469, 2.4941412, -0.8509856, -0.7150132, 1.1363107, 0.8420556, 0.5165584, 0.9273428, -0.0471595, 1.4680234, -0.3598955, -0.4616825, 1.0248003, 0.3652015, -0.6573590, 1.0582744, 2.5048522, -1.4967100, -2.2298935, 0.5501792, -0.4202360, 2.0827222, 0.6689090, -2.3789704, -0.6287612, -1.2052949, -0.6010431, -0.8035681, 0.6742244, 2.6026929, 0.1973211, 2.4146332, -0.1898319, -0.0113841, 1.6744030, -0.3538982, -0.4762931, 0.1315120, -2.0324618, -2.7379363, -2.9679894, 2.4099571, 1.9378028, 0.8737614, 2.1185120, -1.6437462, 0.6222298, -0.5947414, 0.7896893, 0.1706528, 1.5765086, -0.4532455, -2.8757374, -0.0587888, -0.2307883, -0.6978181, 2.1290292, 1.8596632, 2.8950693, -1.0907340, -1.4421818, 1.7264222, 2.3183740, 1.7783099, -1.7014476, -1.9515102, 1.0728816, -0.1855177, 1.1487484, 2.0428653, 1.0315159, -1.5413043, -0.2016704, -2.6750500, -1.2966713, 2.8623806, 1.4365384, 0.2549831, 1.4855898, -2.0660395, -1.4483853, -2.7476584, -1.0270182, -1.3871584, 1.6218063, -0.5313644, -0.5231982, 1.9935972, -2.7062091, -1.1278360, -0.4711964, 1.5320134, 0.7584139, -1.2909608, 1.8808261, 2.8656718, 2.9039806, -1.6750791, 2.9612705, -2.3805690, 2.5434136, -1.3962860, -0.0617304, 0.4651853, -1.3749595, -1.0075677, 0.4506794, 1.9791880, 1.8074217, -2.6489824, 0.2635947, -2.2203723, -1.7650424, 2.8475498, -1.7619474, -2.0352424, 2.2634605, -2.4325465, -0.7366166, 2.7009324, -1.1434817, -1.6013794, -2.7561004, 0.9309827, 0.2654651, -1.7240004, 1.2717805, -0.6925160, 2.2729740, -1.6001293, -1.2693369, -2.6395516, 1.2550150, 2.8766611, -2.2801706, -1.8800009, 1.2400316, -2.2635562, 2.2719376, 2.6542249, -2.6044658, 0.4736363, 1.2891118, -0.2291769, -0.9256012, -2.2185039, 2.9364514, -2.3344481, 0.2333174, 0.9105005, -2.7099949, 1.7621319, -1.4311153, -1.2390335, -2.5942679, 2.5182540, 0.7777382, -2.4284153, 2.9761080, -0.8713521, 1.3591293, -2.8700334, -2.1943570, 1.4916302, 1.9049323, 0.4743409, -2.2803040, 2.3522470, 1.2155226, 0.7212265, 1.5731350, -1.8532370, 0.4155896, 2.1370112, 2.2452721, 0.5617317, -1.1936745, -0.3627916, 0.2775345, 2.9062561, 1.4344766, 2.6675138, -1.9424487, 1.2002495, -2.9008784, 0.0977738, 0.2471161, 0.5155265, -1.0595840, -2.0443857, -1.1381691, 2.4006490, 1.6399939, -1.9280920, -0.8791031, 2.1696531, 0.2242812, -2.9552941, 0.0364486, 2.0267253, -2.7411654, -1.7723511, -1.9255820, -1.7439660, 0.1175864, -0.2144965, 0.9269728, 2.3985230, -1.8553728, 2.1239145, -1.6207289, -1.3359105, 0.5314275, 0.2435965, -0.5521098, -1.3516575, -0.7006594, 2.3509066, 0.1398119, -1.5303737, -2.7710992, -1.4353298, -1.1293456, 2.9476169, -2.3859328, 2.7075688, -1.8753846, 2.5848783, -0.4071647, 0.0875887, -2.7720768, 0.4510331, 1.6450582, -0.8005939, 1.0475492, -0.9210511, -2.9834091, -2.2219448, -1.6231634, 1.2374307, -1.5917716, -0.3021189, -2.0933004, 0.4357954, -2.8572844, -0.4712855, 0.0702012, 0.1689460, 1.5792898, 0.0805712, 1.8920668, -2.1062000, 2.5593154, 0.9228538, 1.8748984, -0.0590776, -1.6850380, -2.7755581, 2.6437266, -2.4161357, -0.2883141, -2.8022082, -1.3716010, 0.2513970, 0.4125490, -1.4821543, 0.7091653, 1.1785113, -0.0927478, -2.9644636, 1.4099555, -2.0455850, 2.0028131, -1.1190274, 0.2352522, 0.1656579, -1.6721151, -2.9060497, -0.4847467, 0.3752808, 1.6075013, -1.2686400, 1.0482117, -1.1836350, 0.0479742, -0.8454985, 1.6162599, -0.9265941, -0.7325993, 1.5278237, 2.6805266, 1.2414188, -1.2350332, 0.5131305, 2.1850545, -2.6223224, -1.2368809, -1.4270044, 2.8522510, -2.3364202, -2.6650321, -1.5233502, -1.3463121, -1.9018724, 0.5153932, 1.3713204, 2.7295490, 2.1957703, -2.5891404, 0.0218758, -2.0782754, -1.5266380, -2.5281897, 1.7130652, 0.4654105, 1.7760062, -1.9079337, 2.9996242, 1.3629968, 1.9940087, 2.3743926, 1.9928644, -0.9036622, -2.8068324, 0.0435246, 0.5079907, 1.7018971, -0.5046101, 2.1955350, -0.8427398, -2.7709563, -2.5957555, 2.5471359, 0.8127968, 1.3116966, -0.5674552, -1.9000132, -0.1851124, 2.5676561, -1.8006851, -1.8944485, -2.1226097, 1.4315911, -2.5930006, 2.8008942, -2.3457920, -0.7118173, 0.5251725, 2.0405298, -1.5866652, -1.1554585, -0.4505501, -2.3673304, -2.9143794, 2.6031522, -1.1682305, 1.0199669, 2.2121614, 2.1875919, -1.7816441, 1.7174965, 0.1022348, -0.1207404, 0.6194139, -1.2140946, 2.2283628, 0.6916288, 2.1768555, 0.7151004, -2.1185866, -2.3022969, 0.1663899, -2.3098567, -0.3176141, 2.2475776, -2.8124884, -1.2806421, -2.5163694, 2.9027011, -0.7728337, -0.7918082, 0.3447607, 0.6416177, -2.6316254, -1.5080775, -0.9998149, -0.7404517, -1.5570948, -2.7378422, -2.6112701, -0.9501830, -1.6797719, -2.4624082, 1.3993827, -0.2678290, -1.7487429, 1.5899409, -1.7254248, 0.7442402, -1.9277707, -2.0504834, -2.1794433, -2.4926998, 1.5180736, -0.5268383, 0.9403541, -1.8014404, -2.6945261, 2.3597757, 2.0116778, 2.0314166, 0.1922273, 2.6446125, 0.4508918, 1.2170551, 0.0771092, -0.0001052, -0.3432194, -1.4530341, 2.8570991, -0.6689875, -2.9214860, 2.4174008, 0.7869963, 1.9455409, 0.6212125, 0.3972611, 0.9423315, -0.3783330, 0.1246163, -2.5273742, 0.6656592, 2.4819860, -0.1797754, -2.7567732, -1.3853656, 2.9359405, 1.3229816, 1.5185875, -1.1205597, -0.9886835, -2.9371216, 2.4914560, -2.5002189, -0.7984874, 0.5688176, 2.1519165, 0.6831796, -1.5021255, -1.1310269, -1.4699343, -2.6251182, -2.6123044, 1.6864335, -0.7603339, 1.5856808, 0.0705816, -1.0142986, -0.8706608, 2.9627512, 0.5987959, -2.4991425, 2.9487570, -2.3827709, 2.2104114, 2.6556818, -2.5351497, -0.7622708, 1.8971633, 2.9960364, -1.3086274, -1.8683965, 1.8696232, -2.6518953, -0.3691668, -2.0686535, -1.6414014, 0.6479027, -0.6355956, 0.1249204, -0.2068156, -0.6897017, -2.4010307, 2.9955168, -2.4279071, 2.1058705, -2.0712869, 0.9946624, 0.8838525, 2.8929842, -2.8992812, -1.0257991, 0.4801837, -2.1224773, -1.6033478, -0.3231856, -2.9104100, -0.5370935, 0.9064667, -0.4366234, 1.7333203, -0.4400962, -2.6102477, -2.8539552, 1.6462525, -2.3818578, -2.2328957, -2.9647050, 1.2378074, 2.1418483, -0.9049962, -2.2235809, 0.1867423, 2.2318304, 2.6389679, 1.3354499, -2.3342738, -2.8316659, 2.4171940, 0.6448082, 2.5724050, -0.9273203, -1.7043836, 0.2269329, 1.9422247, -2.3089002, -1.2469214, -1.5127234, 0.5333913, -2.0547991, 0.4666491, -1.4666607, 0.4733219, -2.1049967, 0.2465934, 0.7995355, -2.8535554, 1.0940852, -1.5786309, -0.2957134, -0.8625288, 0.5056562, -0.9233278, 1.2605035, 1.3765233, 1.5762939, 0.9231870, 1.7270487, 1.0341373, 0.8306855, 0.2079995, -1.0140999, 1.3073603, 1.8900328, -0.7869011, -1.2442346, -2.6851738, 1.0578434, 1.9128451, -1.7401435, -1.8720615, 2.1079523, 2.9475255, 1.8118425, 2.8648128, -2.6867888, 2.2238141, 1.5898076, 2.2852507, 0.3208582, -2.6955270, 0.3321850, -0.5548420, -2.9679401, -0.7769618, -2.4956168, -1.4281428, 0.7008559, -1.1937555, 0.4144542, 1.0956855, -2.6891698, -1.9910970, -2.3994985, -0.1593170, -0.0732109, 1.7811424, 2.3347733, -2.3028159, -2.0996277, -0.1305491, 0.8975162, -1.5957147, 0.9179473, -1.2777235, 1.9987845, -1.8653641, 2.9496869, -1.7520914, 1.0830626, -0.4882887, 2.7776165, -0.5047454, -1.6355546, 1.4354943, -1.9992185, 2.8890025, -2.3404498, -1.6918539, 0.6839247, 1.6014679, 2.1591886, -2.4970453, -0.2896972, 1.9892370, -2.7484664, -0.4614146, 1.6045531, -2.7035992, -2.1027802, -0.4521793, 0.6448915, -2.9221238, 1.8825385, 2.4185272, 0.0461787, 0.6420341, 1.0013410, 1.6283605, 1.9320759, 2.8330514, 0.5606045, 0.4977335, -1.6164244, -2.4887874, -1.1054023, -1.3571558, -2.2219856, -1.9971512, -2.8073975, 1.1442981, -0.3233502, -0.8094399, 0.7473236, 2.3225462, -0.3719873, 1.0151104, 1.0831274, -2.0265506, 1.2501211, 1.3060398, -2.8443047, 1.9809829, -2.0629289, -1.8441711, -0.1369873, 1.5265123, -2.1785970, -2.6375236, 2.2622032, -0.7881081, 1.6332878, 2.8616101, -1.5788488, 2.8164505, 0.2307350, 2.7369268, -0.0163087, 1.2564322, 2.1984853, -0.6201033, 2.3092705, -0.0438906, -0.8357183, -2.2944671, 1.2802718, -0.3178405, -0.2642538, 1.3448767, -2.5035239, 0.9727360, -2.8650511, 2.4868972, -1.8503977, 1.8000899, -1.5321654, -2.1006094, -1.0653625, 0.6141204, 2.7479219, 0.7586992, -0.1709171, -2.1582249, -1.6089671, -0.9464444, -1.9727618, -0.5433165, 0.8902834, 1.0547254, -0.8710257, 1.9105915, -1.4928586, -2.9964013, -0.9213182, 2.7975609, -1.1724690, -1.9262954, 0.7714354, -0.5965328, -2.5918724, -0.5987565, -0.8172008, -2.6908237, -2.0901927, -0.9148383, 0.1441493, 0.3230048, 1.0298149, 2.7542073, -2.3508221, 2.3475687, 1.3420902, -1.3917353, -0.3417977, -1.4610100, -1.5497548, -1.3943047, 2.0370058, 1.0074616, -2.1579881, -1.5456021, 0.1511564, 0.7321903, 1.2039538, 0.7837681, -0.1596375, -2.8667761, 2.7519653, 2.4077737, 2.5658503, -2.7773506, -2.4426046, -2.6023073, 2.3601100, 2.0212081, -1.9366276, 1.3102790, -0.0601227, -2.0315844, 0.9824644, -1.9836385, -0.8179719, 1.9329119, 1.7434081, 1.6239516, -1.4601079, -0.1018544, 2.5770125, -1.1355071, 1.9665431, 2.2716849, 1.4583696, 2.6154844, 1.4127391, -0.1994761, -2.2737283, -1.8050599, -1.1497360, -2.5128759, 1.4010869, 2.8177353, 0.3686645, 1.7379529, 2.1492250, -1.0176242, 0.9780902, 1.2033706, 2.1520158, 1.3101830, -1.0530589, 1.9610048, 1.2897148, 1.0347014, -1.2838516, 1.7637244, -2.1958199, 0.9312682, -0.2576398, -2.9732437, 2.4219710, -0.2540377, 2.4758403, -1.8964497, 0.5064504, 0.0385075, -2.3648159, 0.9208891, -0.9082790, -2.8871790, 0.1590001, -2.8533379, -2.3972125, -1.9188394, 0.3737808, -1.1011445, -1.9416702, 2.7362216, 0.2894375, -2.8484136, 1.3402946, 0.1586861, 0.4369827, -1.1615783, 1.4497000, -0.7740511, 0.9842769, 1.9598966, -1.4505918, -0.3717547, 1.3483063, -1.7046113, -2.8990067, 0.0391238, 0.6816848, -2.1066257, 2.3797904, -2.9394353, 2.9156095, 0.5503899, -2.5519776, -0.0610915, 1.8137740, -0.6731171, -0.1143310, -0.5201018, 2.1592173, -0.1130391, -2.9757706, -0.8961055, 1.2132421, 0.0688717, -0.0373179, -0.0578876, -2.8821004, -1.8828046, -1.5251077, -1.6100947, 2.3883447, 0.6555028, -2.5416228, -0.9546832, 2.0369288, -0.2056974, -0.3952572, -1.4118652, -2.5168543, 2.8885103, 2.0248460, 2.8465269, 2.2701947, -1.0369396, 0.3581585, -2.8501403, -1.8542824, 2.4801660, -2.8350772, -2.6992818, -2.1836601, -0.9294226, -1.1807869, -0.5090387, 1.9510798, 0.1417350, -1.9361113, -1.2795503, 0.9323874, -2.5779156, -1.8701965, -0.6809769, 1.7963537, 0.9559042, 1.1430321, -0.9799620, 1.5513971, -2.5333104, 1.4142928, -0.7735197, -1.5951411, 2.0886508, -0.7951376, 0.8363480, 1.4238062, 0.2424525, 0.6482268, 0.3328889, -2.0113768, 0.5177551, -0.3120138, 1.2259028, -0.2371811, -1.9574060, 0.0262221, -2.9426637, -2.0668412, 0.9702335, -2.6246043, 2.3467070, 1.6726229, 0.0452299, -0.0294553, -0.1616218, -2.1549788, -0.4304100, -1.6092083, -1.2767642, 0.8761441, -1.4855181, -2.2878976, 1.8746110, 2.6370818, -2.9957129, 0.5911985, 1.2635666, 2.5016799, 0.9182172, -0.1308071, -0.8101863, 1.5586916, -0.5154538, 0.5413745, 2.4634671, -1.5139095, -1.9077180, -0.3655919, 1.4711323, -2.3087694, 2.0708535, 2.8918433, -2.1303818, 1.6364812, 2.1292474, 0.7354079, 1.2346364, 1.7485358, -2.4033978, 0.5345437, 0.2221562, -2.9118466, 2.9809127, 2.0113368, -1.7466471, 2.1291322, 2.6764750, -2.8238887, -1.8131562, -0.1313096, 2.7643044, -1.3758553, -1.0913998, 1.4069144, 1.9055488, -2.3967527, 1.9966571, 2.0717398, 2.7415731, -0.5790399, 2.8881973, 0.7693516, 2.5984020, 0.4025558, 1.6662105, -1.0226824, -0.5409758, 0.5488245, -0.4373748, -2.8555587, -0.6781699, -1.3601572, -1.2308146, -0.4926607, 1.2788643, 1.2113755, 2.6030644, 2.6355657, -1.9312571, -2.7716720, 1.0369267, -2.9966973, 2.9291985, -1.8128154, 1.9439993, 2.5845315, -0.8173141, 1.3454034, 2.7813160, 0.1090033, 2.8436046, -0.6176908, -1.6919948, 2.4757179, 0.7495127, 1.4149414, 2.5479256, 0.5777931, 1.1401899, -2.2506790, 2.0118083, 1.4331485, 1.1340709, -1.7801880, -2.5288548, 0.7472129, -2.4140647, -2.4334488, 2.1156802, 0.4369620, -0.8646029, 2.9159973, -1.7775685, -1.3708763, -1.0956992, -0.0862207, 1.4183029, -0.3318820, -1.4746751, 0.1013437, 2.1319846, 2.0358290, -2.9279829, -2.7950666, 0.1176947, -2.2214576, 1.8807300, 1.3665706, -2.3361326, -1.3846711, 1.2389083, -0.1972800, -0.0740040, -2.9543065, 0.8309665, 1.9315870, 1.2448543, 1.0660523, 0.9136173, -0.3663817, 0.3010993, 2.3263550, -2.9000408, -0.2888338, 2.9215108, -2.5885480, 0.7833677, 0.8042193, 0.4411333, 1.5469714, -0.1361784, -0.5448018, 0.0105709, -2.0448236, -1.0344612, -0.0406012, -2.2963123, -2.7503815, 2.9549003, 0.7310315, -1.6897184, -2.7093517, 0.7574172, -0.7846213, 0.1329291, 1.5509599, -2.2516368, 1.4805239, 2.5769930, 2.9258806, 0.1503613, 0.2020983, -1.4294170, 1.5867595, -2.3747433, -0.6787509, -1.3009289, 0.8831771, -2.0483096, 1.7227370, 1.8237018, 2.1443821, 2.3450866, -0.5569588, -0.7708829, 1.7835676, 1.3215308, -0.4672171, 0.9921298, 1.5451640, -0.9318341, 1.0625554, 1.9728096, -2.5442181, -2.8029202, -2.7083536, -0.4143666, -1.7619748, 0.1595520, 0.4263924, -0.2280029, 1.9742660, 1.5126153, -2.7547769, 0.9550488, -2.5175924, 2.8487830, -1.5541046, -1.8393710, 2.9786229, 0.5383529, -0.1045984, 1.5639867, -0.4961050, 2.4987477, -2.9507101, -0.3217799, -0.9671033, 2.4761067, 1.2846669, 1.5686852, -0.0451190, 2.8507023, 2.2465744, 0.0960458, -0.3422782, -2.6399065, 1.1488104, -1.9893708, 2.8325947, 2.0996987, 2.5730623, -2.2365776, 1.8264543, 2.7073191, -2.5542015, 2.9844654, 2.1372757, 2.8926952, 1.3662627, -1.7918496, 0.6352801, -0.6494549, 2.1813146, 2.2354700, -0.1847703, -1.0070440, -0.1661446, -1.7660103, 1.0869868, -2.9703352, 2.0908290, 1.9606207, 1.2018781, 0.5559215, 0.2752661, 0.9097975, -0.6667126, 1.7113018, -2.7620174, -2.0020509, 1.0969889, 0.6360870, 2.2304028, -0.0792432, -0.7929124, -0.1945227, 1.7280729, 1.4872908, 0.6964357, -2.8362543, 1.0870926, -1.9689065, -2.2615907, 2.8337123, 0.9140677, 0.4806942, -2.5222158, 2.6206580, -2.9037886, -2.2551768, -1.1530109, 2.8533057, 0.0669418, -1.7797672, -2.3479241, 2.2707234, 2.1055198, -1.0443203, -2.9834850, 0.8498336, 1.7119014, 0.3118453, 0.4536055, -2.7839810, -2.4988018, 2.8608845, 1.4881320, 1.5108971, -1.9240174, 0.0473251, 1.9757212, -2.8535383, -1.8366029, 0.4515891, -0.4342518, -2.2808318, -1.6909818, -2.5468052, 1.1939632, 0.4181058, 0.0454793, 2.4161613, 1.4610656, 1.2699167, 2.4106481, 0.4538850, 2.9159128, -0.9418628, -2.5965465, 2.5094289, 0.3347516, 1.8884935, 1.6837711, -0.3113533, 0.6710531, -1.9289382, 1.2977667, 1.1687435, -2.6660815, 0.6743330, 2.9151650, -0.5266356, 0.9675795, -0.6191047, -1.0231272, -1.8578409, 2.2954454, 0.6954182, -2.8973859, -2.6638238, -0.1574303, -0.4671948, 2.3753673, 2.8857303, -1.8854305, -2.5439708, 1.4682003, -2.0031017, 2.8133287, 0.9414684, 2.9722093, -0.7674627, 2.6598360, 2.3238362, -0.4562033, 2.7142865, 2.1696487, -2.7630661, -1.6302001, 0.1876428, -0.9603304, -2.2550125, 1.8451406, 1.8673377, -1.9104779, -2.4866331, 2.4443497, -0.6931715, -1.3228692, -0.3528999, -2.7696338, 0.4011820, 0.6960817, 1.6468364, 0.9827314, 1.4132176, 1.2084813, -1.1599808, 2.0169194, 1.4849186, -1.7097704, -2.2639837, 2.2462441, -1.2053269, -0.2619170, 1.4758350, 1.1052060, -0.4636770, 2.1846508, -1.3458278, 1.9309286, -1.3776128, -2.3177669, 1.5471388, -2.1077578, -2.1209643, 0.7556955, -0.7734798, 0.3915237, 1.9429830, -2.7439223, -1.4864263, -0.8985790, -1.0421177, 2.3474955, -2.9698352, 1.4148753, 1.3285241, -0.1221131, -1.9562762, 0.7998601, 1.2527407, 1.4575730, 2.1688493, -0.3978770, 1.8476728, -0.9142573, -0.0659087, -0.6734391, 2.0376214, -1.5709749, 2.5632085, -0.7245312, -1.5620004, 2.1681478, 1.8081103, -0.9160850, -1.7638398, -1.1783379, -2.7179699, -0.0745100, -0.0058204, 2.3868326, -1.1528762, 1.1677633, 2.0728654, -2.7726550, 2.8526143, 2.2131791, -0.4124675, 2.1354960, 0.6346587, -1.6089134, -0.7072617, 0.1677383, -0.9620335, -2.5237011, -0.2600416, 2.0233000, 2.4339858, 0.5404053, -0.6801051, -0.0180003, -2.4670422, -2.0319807, 2.4127209, -2.5710265, -0.7851545, -0.1399026, -2.3556701, 0.3900230, 2.1332541, 2.2546682, -0.3703302, -0.4193346, 1.2375995, -0.2971422, -0.6820948, -1.0533596, -1.4814538, 1.4947716, 1.8390019, -2.0300051, -2.4421302, 0.3335079, -1.2558865, -1.4892685, 0.1546982, -0.1522429, 0.6018952, -0.1762999, 1.8130906, 0.8770100, -2.7891660, 2.0616558, 1.9232655, -1.4736716, -0.7412949, 2.3641035, 2.9826960, 2.8645223, 2.3146490, 0.5943730, 2.1611770, -0.2325000, 1.2223678, 0.1605285, 2.1912174, -2.6827932, 2.7761738, 0.5582975, 0.2286272, -1.7736854, -1.4486357, 1.9082113, 1.9629369, -1.5411824, -1.6323406, 0.8166739, -2.6301056, -1.3127206, -0.9806812, -1.5400010, 0.3307035, 0.6748367, 1.8825910, -1.8452041, -0.6745623, 2.3877597, -1.1677917, 0.7889368, 0.1976767, 2.5967404, -0.0538178, -0.0520211, -1.3499057, -1.6415599, -0.3131987, 0.7484665, -0.3778768, 2.1841381, -1.1020955, -2.7409598, -1.7288042, 1.8987346, -2.4863215, 2.4357245, 0.7956468, 2.5438516, -1.3079952, -0.8993368, 0.2363495, -2.6806283, -2.7867839, -0.2140291, 0.8666689, 2.9009738, 0.9075391, -1.3445071, -1.6853342, -1.0333592, -2.4992488, 0.6691530, -0.1668068, -2.6232398, -2.7414884, 0.0992035, -1.7809740, -0.3927308, -1.5496116, 0.8702048, 2.4811197, -0.3153418, 2.8038004, -1.1559628, -2.5831251, 0.2481634, 0.0467305, -2.7590624, -1.3651349, 0.1681989, -0.6017435, 2.2970051, 0.9527078, 2.6036937, -2.5014657, -2.0029883, -0.2388975, 0.1698165, -0.4580450, -1.1086744, -0.9785804, 1.4227326, -2.7262278, -1.1157781, -0.8644691, -2.6585492, 1.8852454, 0.0343922, 1.2146712, -2.2878308, -0.9333150, -2.7695616, -1.3796358, 0.2408932, 0.2888706, -0.0130725, 2.1918604, 2.3958402, -2.5281453, 2.2405481, 2.3323479, 1.0671860, 2.1312561, 2.4196840, -1.1903047, 1.2361034, 0.1656145, -0.0085500, 2.4023889, 1.5734369, 0.7340043, -1.3902368, -2.9932397, 1.8370332, 2.5024932, -0.5914956, 0.4045236, 2.1192079, 2.7033275, 1.6997719, -1.6714356, 0.2000449, 2.3481788, 1.6592237, -0.4866147, 1.6885220, 2.5068104, 1.2285026, 1.5452455, 2.8442832, -2.1245728, -0.8157842, 1.6505506, -0.8402851, -0.2157801, -0.7900673, -0.3560318, -0.7543018, 2.2183696, 0.8411889, -1.3208736, 0.8179255, 1.6361116, -0.1948057, 1.9786219, 0.2604136, 0.8019765, 2.2821698, 2.5042836, -0.1491440, -2.6889393, -1.1735454, -0.3821551, -0.4637076, -0.9625552, 2.1661600, -2.5101825, 1.7047486, 0.8399195, 1.8518348, 2.4475912, -2.4212530, -2.2085230, 1.7560975, 2.6625157, 2.1443047, -0.6261913, -1.2738391, -2.4889994, 1.2875457, -1.9859470, -2.9994150, 1.8854128, -1.3646463, -2.6694979, -1.6697832, 1.5363429, 2.5733597, 2.5016698, 0.0941535, -2.6255413, -1.1936073, 1.1978686, 2.6036801, -0.2025330, -0.4192153, 0.6616185, -1.4173158, 2.5379892, 1.2305375, -1.1731079, 1.8376804, 2.2389073, -0.8479233, 1.5840280, 1.0844075, 0.8536962, -0.1944611, 2.1933093, -2.0523333, -0.0152400, -2.8324101, 2.0180151, 1.9198416, -2.8680436, 1.9122353, 2.9012396, 1.4938326, -0.3940943, 2.5667870, -1.8256468, 1.4659953, 0.9841919, 2.3766003, 1.6183564, 0.0309956, -1.0555142, 2.9649243, 2.3122259, 2.5877357, 0.1910901, 1.9315656, -1.7425738, -0.9101854, 0.0591621, 0.5954963, 1.2038455, 2.3219669, 2.4756347, 0.4303245, -2.1638678, -0.6354044, -2.8745810, -0.8229687, -1.9569482, 2.3463656, -1.6328573, 0.9588202, 1.6150647, 1.1207473, 2.4168720, 2.5869463, 1.9670530, 0.5748116, -2.2856139, -1.0137052, -2.2155228, 2.7263096, -1.1288885, 2.1583608, 0.7484514, -1.6915519, -2.2546611, 2.0143754, -2.9914381, -1.9287530, 0.6262276, 0.6638558, -2.2076173, -1.2112313, -0.4889581, -1.6063519, 2.0300889, -0.3112100, 1.8244294, 0.5871901, 1.3481544, 2.1629360, -2.3949131, 0.6500102, 0.9410756, 2.5217466, 0.6267721, 0.9477030, 1.6461950, -2.8318787, 1.6169749, 2.2279761, 1.4599431, -0.8331887, -0.5625409, -0.0684263, 1.4950046, -2.7851652, 0.1770234, -2.2966968, 2.4602331, 1.5446016, -2.4650385, -2.2033630, -1.8307990, -2.4747701, 2.4061504, -1.0609164, 0.1042248, 0.8674757, 0.7691920, 2.5264431, 2.1542468, -1.8448012, 1.6347857, 0.1412949, -0.4915612, -0.2797668, -2.5956494, 2.1406781, 2.9327442, -2.1291079, 0.0135658, -1.0951113, 0.6379483, 2.7275992, 1.0875355, 0.9509770, 0.0692550, -0.9196259, -0.4682032, -0.6120989, -2.6420078, -1.8278171, -1.5934974, 0.4333696, 2.3588175, -0.0285681, -1.2965414, -2.3961805, 1.7216577, 1.5074370, -2.4812857, -2.1407760, -1.4377784, -1.1986198, -2.8901550, 0.7063575, 2.6098435, -0.7845635, -2.1498543, 0.0925009, -0.7176131, 1.3864291, 2.1518998, 1.9302673, -1.5659990, 0.4800525, 0.2410215, -0.9128529, -2.7523346, -2.2133208, 2.4779471, -1.1607443, 1.9827940, 1.4723452, 0.4460924, -2.3131434, -0.7677749, -1.0434246, 2.9324696, 1.1903504, -2.7113102, 1.2564115, -0.0511229, 2.4677267, -2.9890894, -1.8440386, -1.6898890, 0.2970270, 2.9451081, -0.2511012, 0.1025319, 1.4447198, 0.2308670, 1.7688687, 2.4288927, -1.5732153, -2.7513704, -0.3418970, -2.5495958, -0.6064139, -1.3379757, -1.4722160, 1.4059743, 0.0346661, -1.5500241, 1.0952519, 1.3012908, -0.0744523, -2.1165333, -2.6638355, 0.5828283, -1.7790244, -0.2760689, -2.4156356, 0.8548935, -1.6865559, -0.8406061, 0.7965001, -1.9129391, -2.6658138, 2.9107751, -1.1064901, 2.8323635, 1.5445497, -2.0178148, -2.6707820, 2.4504686, 2.4844205, 0.5133783, -2.3082168, -0.3936831, -2.7913923, 2.0574998, -1.9958876, -0.5847310, 2.0046298, -0.7921726, -0.3201773, 1.2521221, 1.7530029, -0.1323006, -0.7475345, -1.0121541, 2.8121481, -0.2621944, -1.3558586, -2.0159486, -0.8625356, -0.1563110, 2.6286757, -2.1775002, -0.9945606, -2.3979525, 0.9349700, -0.3695140, 2.9646741, 1.8434009, -0.2515802, -2.5010935, 1.5225265, -2.3942589, -2.0189659, 0.3560485, -2.0954999, -2.1572863, -0.9972213, -2.8517689, 1.8803052, 1.2388723, 0.9491565, -1.3634795, 2.6019959, 0.0902169, 0.6239821, 1.5440135, -1.1868316, 1.2424328, 0.7400573, -1.5819820, 0.1481055, 0.9373448, 2.6860373, -2.5317938, -1.5286991, 0.6724324, -1.8732673, 0.3817546, 2.5352539, -2.7701910, 0.0848583, 0.0040951, 1.7815798, 1.9633161, -2.7470810, -1.0978169, 1.2583191, 0.3150261, -2.4759509, 2.4438463, 1.4176091, 0.1050439, -0.5243698, -0.5156843, -0.6928085, -1.8134192, 2.3157163, -2.3683979, 0.2212445, 0.1609494, 0.8716249, -0.4416575, -1.6209246, 1.4301042, 1.8806497, -1.6914352, -2.5971244, 1.4954479, 1.1953293, 1.1765975, 1.7829710, -2.3131121, 2.1908525, -2.6233747, 0.2801310, 0.5589546, 2.3896755, 2.3053053, 2.3077977, -0.8515467, 1.1791936, 0.7994432, 0.8063239, 0.3020011, -1.3938206, 2.0922291, -0.3755631, 1.5768413, 2.3083640, 0.7496778, -0.7521404, -2.3639936, -2.3448437, 1.0111342, 2.4914739, -2.3152895, -0.4802523, 2.1419207, 1.9941897, 1.6744409, -0.8527634, 1.0753816, 2.0676878, -0.4717035, -1.0910922, -0.8548061, -2.9086970, -1.1617958, 2.4166287, 0.0577340, 2.1029386, 0.5678418, 1.3974458, -2.0466054, 0.9908447, 1.1033456, -0.2859757, 2.3247342, -2.7612037, -1.4382336, 1.8083410, -0.7557624, -1.0783414, 1.4074706, 2.9740681, -2.1408201, 1.4005553, -0.8558382, 0.0647195, -0.7696295, 0.7971041, -2.5304281, 2.6530570, 0.5919541, -2.9912570, 0.7299087, -2.7103201, -1.7308525, -1.5425726, -0.8220102, -2.3379102, 0.3225150, -1.8192085, -1.2213605, 2.8143252, -0.5986808, 1.3925469, -1.1007177, 1.4290946, -2.6734036, 1.4194941, 2.4208151, 2.3888190, -1.5595129, -1.3938323, 1.0635347, 0.7203230, -0.3020542, 2.0034476, -0.1436585, 1.4711682, 0.5162797, -1.9781791, 1.1795787, 2.9437758, 2.0478943, -2.7711245, 2.8519223, -1.0401271, 2.5348545, -1.7336368, 0.5281288, -0.6177084, -1.0483206, 0.4818500, -0.8144033, -1.4180641, 0.2586095, -0.1825073, -1.3011661, -0.6707540, 0.0284793, 0.7483436, -2.1632311, -2.4681825, -0.7837300, -2.6572904, 2.4841805, -0.1378683, -0.7344512, -2.0907069, -0.7331943, 2.9912435, 0.3778713, 0.7196405, 1.0204413, 0.4185023, 1.2958363, -1.7518565, -1.3615180, 1.8397162, -1.0675615, -0.2244151, 0.3121067, -0.4246800, 0.0489191, 1.2217682, 1.1989235, -2.0009865, -2.0834600, -2.8768180, -0.7265778, -1.9040617, 2.6771482, -2.3121907, -1.5033537, 2.2593710, 0.3927043, -2.0686633, 1.4108256, 0.3349153, -2.5073589, 0.6637675, 0.1708211, -2.8866309, 0.9001250, -0.3539056, 2.5422094, -1.9806870, -0.3082144, 0.3972371, 1.3749771, -0.3625688, -2.1563667, -1.6075328, 2.3010202, 0.9271058, 1.4241965, -0.0733380, -2.4076509, -2.6620055, -0.0974764, 1.3785298, -0.3825348, 0.8333888, 0.6337793, 0.9214063, -0.2811347, 0.0506859, -1.8575255, -1.0225586, -2.0078790, 2.1241802, 0.7104298, 1.0033921, -1.3897291, 2.9794910, 1.7067590, -2.8495945, 0.0993124, 1.3482692, -2.9333585, 0.0709844, 0.5919468, -0.4551418, -0.3608076, 2.6877651, -2.7275537, 2.1629949, 0.1498035, -0.8917360, 0.2563687, -0.3734118, -0.3498961, 0.2961102, -2.7030213, -2.6015885, -0.1568116, 0.0310471, -2.3463047, 1.0064694, -0.9072822, -0.8539527, 1.4552681, 1.0461489, -1.4548403, -1.4044879, 0.2346679, 1.8530252, 0.8064739, 0.5326813, -0.4053247, 0.9615818, -1.9868437, 2.7595112, -0.1894710, 2.4124870, 1.2740233, -0.2228767, -1.9357169, -0.3051083, -2.4554561, 1.4533013, 1.0189192, 0.5250559, -2.0213501, 1.6453094, 0.3250424, -1.9790863, 0.2512605, 0.5364850, 2.4078741, -0.2763177, -1.7359760, 1.7590903, -2.4796818, -0.5090735, -0.4306546, -1.6959775, 1.7891867, 2.1676668, -2.8750338, -0.2972837, -0.2390213, 0.2445069, -1.6237136, -2.1962311, 0.1378258, 2.6677849, 2.0728053, 0.0692706, 1.7733688, -1.7069823, -0.5677632, -0.4361161, -2.4422457, -0.9558275, -1.6943249, -0.0150526, 1.7738876, 0.3027963, -2.4643884, 2.0120411, -1.2532941, -1.8842287, 0.0437886, -1.4794456, 0.5412934, -0.2186091, 0.8740193, 0.7637330, 2.5288967, -1.4911117, -2.0530548, -2.0061277, 1.0429037, -2.8405530, -1.1155971, -2.2757761, -1.3781830, -0.5156362, 1.6197025, -2.8879231, -2.8017846, -1.1437705, -2.1233923, 2.6091453, -2.2529504, -1.5545757, -1.7419797, -1.7787483, 0.8349384, 2.7154859, -2.5632368, 2.1898237, 0.5598518, -0.9645701, 2.7305696, 0.7422308, 1.7415272, 1.8440542, 2.5941789, -0.1743683, 1.8624211, 0.7139842, -1.7974145, -2.3180347, -2.7593374, 1.8848039, -2.1087549, 1.3458120, -0.9341667, 2.4019866, 1.6210471, -2.7734754, 0.2779727, 1.2721007, 2.5311925, 0.4287928, -0.5887688, 2.2764722, -1.7309167, -2.7277358, -1.3905016, 0.2250527, -1.1677538, 1.2824890, -1.2707790, 2.4328910, 1.8178993, 1.7289215, 1.7735417, -1.0438863, 0.0721965, 2.1040256, 1.6484373, -1.8647890, -2.6381304, 0.4250465, 0.1605380, -0.1778200, 2.6645445, -0.7087222, -0.6470688, 1.7080352, -1.7021435, 0.9877663, 1.7760033, -1.8887270, 0.4173496, 2.5376349, 1.1098126, -1.5972482, -0.2550238, -1.6182253, -2.6747986, 0.2929087, -1.1233320, 0.4586305, -2.2612966, 2.1570160, -2.5422124, -2.1037301, -1.2184475, 2.9442695, -1.6456689, -2.1674163, -0.3793766, 1.6117894, 0.8708144, 1.1279742, 2.1350804, -0.3298484, 2.8437446, -2.2188276, 0.0209774, 2.8852618, -0.3793233, 1.7353658, -0.0989461, -0.3558092, 2.7999945, -0.5357751, 1.4438234, -2.1723263, -2.5136430, -1.7894173, -0.7981037, 0.1009530, -0.7749156, -2.9092002, -1.7572679, -0.7584830, 2.2031865, -0.1481780, -1.3109979, -1.6673155, 1.0474500, -0.0728512, -0.3519395, -1.7122119, -0.0163723, 2.2512155, -1.6176619, -2.8291417, 0.2736726, -0.9785099, 2.4678372, -0.6613952, 2.7305781, -0.1013191, 2.7884505, -1.5073075, -1.9918302, -0.7350522, 0.3097744, 0.7941621, 2.0015923, 2.0922200, 0.5069873, 0.9708455, 0.3548990, -2.5451872, -0.1241005, -2.0988329, 1.8434701, 0.1253575, -0.6280466, 0.4698549, 2.3251413, -0.7659952, -1.6338202, -0.2615997, 2.3468502, -1.1353449, -2.0737102, 1.0616143, -2.5781463, -0.8864152, 0.1234529, 1.6558132, 0.4364972, -0.4255847, -1.9630523, 1.6106667, 0.5191466, 1.1476844, -2.3491510, -2.6597060, 1.0327095, -2.4623176, 2.4295609, -1.0210541, -1.4044601, 2.0622369, 1.7486590, 1.9170213, -2.5925197, 1.9403657, -2.5670441, 0.9833016, -2.9515912, -0.0579885, -2.7748118, 2.5183934, -1.5327743, 1.5762546, 1.0110896, 1.8588842, -2.8116949, -1.7567798, 1.9239994, 2.1042787, 2.4127223, 2.6899986, 2.5242070, -2.3227597, 1.1849677, 2.2420725, -0.9908857, 1.5545943, 2.7821793, 1.5579635, -0.5279741, -0.7119995, 0.7414159, -0.4823115, 0.6893878, -1.9279273, -0.5699941, 0.2621069, 0.1809981, -2.9097697, 2.4169657, 0.8658306, 0.8619317, -2.9389271, -0.3803068, -0.8590616, -1.6305960, 1.9931474, 1.1515256, 1.7497906, 0.7378704, -2.0457024, -1.7537900, -2.4265192, 2.4741872, 1.0424484, 0.3055177, -0.7826997, 1.9029423, -0.5714680, -2.8499272, -1.6456301, 1.7227285, -2.2208404, -2.5791855, 2.1879044, 1.6513040, -0.8835154, 2.1225944, 0.7977285, -1.2272765, 1.3829158, 1.8224077, -1.7023611, 2.8699087, 2.7054097, 0.4657248, -2.0130238, 2.9859232, 0.8988641, -1.1121438, -1.2524178, -1.5341909, -1.0590878, 1.3585310, 0.6199539, 0.8132450, 2.1425989, -2.1663060, 0.0525765, -2.7176635, -2.4137562, 0.1596648, -2.7872836, -1.8554031, -2.9035096, 2.1219099, -2.8584414, 2.9678101, 2.5853750, 1.0957426, 2.3964253, -1.5497184, -1.6449938, 0.1713289, 2.1262140, -0.1745341, -1.1448509, -0.6339707, 2.5652386, 1.9415026, 0.0241365, -2.1507159, 1.4074274, 1.2383176, 1.4605671, 0.0825146, -2.4933998, -0.6512904, 2.6198319, 0.8782359, 2.4261867, -0.4133875, -0.4365479, -0.1764975, -0.3570678, -2.4815661, 1.5578783, -0.5657697, 1.3717540, 1.8909941, 2.6763595, 0.0986025, -1.9684173, -1.2184900, 2.8529046, 0.1763144, 1.9275569, 0.9597810, -1.5030259, -1.8110949, 0.2511612, -2.7032152, 1.3601779, -1.2096650, 2.1094397, -1.1512239, 2.7746642, -2.9098161, 1.6740444, 1.3244271, 1.0290314, 1.6922917, 2.2109449, 0.3979142, -2.9199508, 2.4437260, 1.4391098, -0.9632288, -1.6907540, 0.1763171, 1.9194523, 0.7134522, -1.3927526, -0.2463056, -1.9343049, -2.4459953, -2.8045050, 0.6763873, -1.4869682, 2.1162378, -0.0105471, -0.8618439, -1.8577176, 0.8376638, 1.6724347, 1.4363137, 0.9696254, 2.9005281, -0.7850788, -1.6328975, 0.7073718, -1.0042369, 0.5347999, 0.2011505, -1.4368940, 2.4793690, 2.3432307, 2.3559324, 2.5130361, 2.6375621, 0.1317601, -2.1567957, -1.1390571, -0.1727770, -2.7765643, -2.2382528, -0.8738810, -2.9370385, -0.6371732, -1.9883444, 0.3260118, -1.6914567, -0.8624834, 2.4649313, -1.7136132, 2.8936905, 0.9882243, -1.1333044, -1.2192865, -1.6461216, -0.2996890, 1.7561181, -2.6302151, -2.8136993, 2.1167101, -2.4105997, 2.1088475, 2.7788477, 1.8398036, -1.1816676, -0.6371225, -1.5684390, 1.8769792, -2.4682022, -2.2431265, -0.5016086, 1.2836591, -0.9990093, 1.5385692, 2.3501452, 0.8615898, 0.7786243, 0.9905267, 0.1604885, -2.4742130, -2.1967567, -1.4529476, 2.3727451, -1.9611224, -2.7353271, -0.2654289, 0.8789446, 1.2195058, -2.0137363, -1.7368303, -0.3325183, 1.7489282, 1.7805879, -0.7986276, 2.1293769, 0.0883985, -1.1091501, 1.8476276, -2.5509299, 0.5151944, -2.4741184, -1.4710052, -2.0524455, 0.8616868, -0.7741196, -0.3412198, 2.9828934, -2.6837039, 0.3342954, 1.2826324, 0.3437817, 2.7503206, -2.8822879, 2.6462335, -0.2043307, 2.6536081, 1.7336501, -2.5485550, -0.4379721, 0.6531441, 1.0473620, -0.3470442, -0.8225420, 2.7648197, -2.4100991, 1.1920446, -2.5255821, -2.9192573, 2.8844306, -0.7710823, -1.0677958, 2.1076720, 1.9466607, -0.0905213, 2.3746267, -1.3628603, -0.5810319, 0.5926830, -2.8906279, 2.0519676, -0.1397037, -0.0029653, -0.0274972, -0.8028946, 1.2965958, 0.6862017, 0.8103730, -2.3796213, -0.5915179, 2.7872950, -0.1817532, 0.0152265, -0.1727835, -0.2330993, 2.7307689, 0.5793135, -2.3416708, 0.6632484, 2.9659347, -0.4464721, 1.6794723, 2.5981358, -2.1733107, 0.1907461, -1.2834083, -0.4165154, -1.5858688, -0.2897749, 0.0286384, 2.3214556, 2.0398355, -1.2341705, 1.5765326, -1.6876658, 0.4841346, -0.4071882, -2.6655335, -0.3909357, -2.5859035, 1.9828299, -2.8949833, 1.9582863, -1.3877110, -0.2574906, -1.2389949, 1.3298369, 0.7924048, -0.8383441, -1.6758418, -0.2585227, 1.2041421, -1.2733079, -2.9527157, -1.5849973, -1.5081653, 0.9919171, -0.9959278, -1.4395926, -1.5325937, 2.2713508, 1.9667143, -1.8276061, -1.2184148, 1.6693284, -0.1023723, -0.4851752, 2.7178118, 0.1012128, -2.7388054, 0.2331535, -1.5356795, 1.0156517, -1.6036219, -1.9331392, -0.5649297, 1.3578239, 2.5498622, -0.0088499, -1.2859091, -0.5321679, -1.0311899, 1.5900532, 1.2414726, 0.3340958, 2.2000296, 2.6122471, 1.7616546, 1.2904890, 0.2487170, -0.8437340, 2.6755261, -1.3343809, 1.7000170, -1.7960261, 0.1383436, 1.0255897, -2.8455875, 1.5047899, -1.8841525, -0.7274294, -1.7692698, 1.5198647, 1.7721781, -1.2084631, -1.0582617, 1.8417686, -2.8610740, 0.1616220, 2.6908265, -1.9185845, 0.7541756, 2.0531194, -2.6610606, 0.0359891, 1.2676030, 1.9697792, 2.0463478, 2.3731938, -2.0665697, 2.9339344, -2.5285980, -2.5894071, 2.6927891, 1.9503023, 2.8657723, 0.3917116, 1.4903580, 0.5716802, -2.6793664, -0.7539681, 0.6164769, -0.2135702, 1.9396859, -2.8155322, 2.8041232, 2.1714780, -1.7430049, -2.9442131, 0.9001797, -0.3076566, -2.7836511, 2.9328289, -1.0981474, 2.8698680, 1.9014319, 2.7189207, -2.5535262, -1.1991717, -1.3486471, -0.0504213, -0.7646888, -2.0607163, 1.0819108, 2.8696742, -1.0505162, 2.9066236, -2.7510350, 1.6478495, 0.5566438, -0.6752135, -1.7054362, -1.8573973, -1.2624659, -0.7264545, 0.1383749, -1.8043015, -1.1083661, -0.2545470, -1.7770100, -1.8551712, -2.7167248, 1.3010857, -0.6057098, -2.2982386, -2.5921243, -0.8018885, -0.4531680, -1.9471667, 2.6131047, -1.1541846, 1.2849274, -2.9344797, 1.6588980, 0.4560499, -2.0595384, -1.5245099, -2.6692217, -0.5263784, -1.4017707, -0.7152988, -2.0925631, 2.1886578, -2.1014979, -1.2954467, -2.0177981, -2.5273821, 0.8100782, -2.9327407, 2.0555462, -0.2160201, 2.3989267, 0.9602900, -2.4203118, -0.9917741, 0.4103010, 1.2890761, -1.6740092, -0.4384980, -1.2940368, -0.2052418, -2.9874651, -0.2700419, 2.7244671, -2.6276437, 2.0016804, -1.1293988, 1.3312225, 1.0510419, 0.0995523, -0.5359634, -1.2072785, 2.8564610, -2.6724308, -1.1277544, 0.7680411, 2.6205371, -0.7728516, 2.7929209, 0.4329117, 0.7535563, 0.7316461, 1.6190068, 1.6105907, 1.0879688, -2.8938933, -0.4491507, 1.1267694, -1.4284414, -2.0810697, 1.4882515, -1.1651023, 0.5469824, 1.3469362, -0.1370003, -2.1060769, 1.5836804, 2.3288432, 1.7263416, 1.7876840, -1.8543815, 2.8969202, -0.4828994, -1.1876791, -1.4632113, -1.2245548, -2.6243865, 1.9357231, 2.0436147, 1.8553386, 2.1675509, -1.5152192, 0.9261860, 0.3115984, -1.3752832, -2.2617353, 0.4940693, -0.9700721, -1.4598806, 1.1941241, 0.4984214, -2.4010161, 1.6008480, 2.8841035, 0.5086707, 1.6884063, -1.1712323, -2.1502802, -2.8394908, 1.3302750, 0.6290208, -2.1937596, -1.3638986, -2.2475611, -2.7472627, -1.0097721, -0.2022422, -2.7679346, 2.5063368, 0.5264328, -2.6299330, -0.2187940, 1.5144490, -1.2421673, 2.6941339, 0.4807515, -0.1049229, 1.2227600, 2.4161441, 1.1862377, -1.0418889, -1.4209955, 1.0409180, -0.3800605, 2.5077852, 2.1292573, 2.9031181, -2.5898065, -2.2183184, 2.1134321, 2.3010471, -1.5981047, 2.4784698, 1.0276178, -2.0633594, 2.6252880, -1.1722038, -2.1378993, 2.0560588, -0.5581800, -0.7811252, -1.7541068, 0.3629659, -0.7723031, -0.0746687, -0.8340444, -1.3117619, 1.0817788, 0.2808188, -2.5728571, -1.2580149, 1.1062866, -2.8740353, 0.5712372, -0.8330685, 0.4244640, -0.8475219, 2.1116304, -1.3326628, -1.5147629, 1.1360684, 0.3684525, -0.4757214, 1.2695235, -1.1102357, 2.2636935, 1.6837667, 1.0142641, -0.3413419, -2.1040259, -1.0557358, 2.5555817, -0.5544193, 0.0407008, -1.8998583, 0.6630994, 2.3625384, -1.1066079, -1.3792263, 0.9764388, 0.5220176, -0.1848629, 1.3151776, 2.9558203, -1.1531776, -0.0570252, -0.1890265, 2.7410013, 0.6573516, 0.6034930, -2.1751149, 1.6181991, -0.0075982, -2.0580716, 0.6567017, 1.8476249, -0.4753415, 0.1758645, 1.8296680, 0.7695571, -2.1140589, -0.3658746, -2.2986659, -1.3261037, -0.9692397, -2.2144154, 2.9700182, -2.4781427, 1.5086239, 2.6270797, -1.3838204, 1.3752036, 0.5399959, -0.2724070, -0.4041802, -1.8603515, 2.3028472, -1.4429385, 0.4457534, 1.5608837, 1.6765379, -0.5986676, -1.0414010, 1.3530894, -2.9507800, 2.6404983, -2.2964419, -2.1531782, 0.0045617, 1.0337917, -0.7395752, 2.1129221, 1.3046300, 0.1740726, -2.7411503, 0.1804607, 2.3297938, 1.1446513, -2.3607939, -0.3262464, 2.1720934, 0.2866483, 2.6781201, 1.4843186, -2.4161745, 2.4675397, -0.2923528, -2.4081907, 2.4770644, -1.4330900, 2.2670931, 2.8428323, -2.3539128, 0.6354678, -2.7178591, 1.1453256, 2.6674121, -1.4994080, -2.6342788, 0.1139780, 0.9153643, 1.4853145, 1.7206667, 1.9113023, -1.4391331, -0.5791746, -1.0311759, 1.6893142, 2.2574190, 2.6601791, -0.6780811, -0.1818913, -2.2603332, 0.1004326, 2.5912104, -1.1034103, -0.0684234, 2.4405303, -2.9399860, 0.0299332, -0.6242184, 0.6523300, 2.8851821, -1.9764807, -2.1337022, -0.8880521, 0.2040520, 2.5402721, 2.3567564, -0.2872788, -1.1584435, 1.3319196, -0.1556526, -2.3520036, 1.0411490, -2.3740079, 0.8519936, -2.3559724, 0.4295736, 0.0240250, -1.1152819, -0.7182048, -0.9042871, -0.3013077, 1.8333316, 1.4401734, 2.4308445, 1.5806517, 0.0829045, 1.4284816, 2.3687919, 1.5928663, 1.8702273, 0.4200304, -2.9094423, 1.0175222, -2.4652166, -0.2335365, 1.4298778, 1.3187241, -2.3454720, 1.8649719, 1.3012424, -2.8029675, 2.0442222, 1.6594542, 0.6028346, -1.6615853, 0.2324484, -1.2141894, -0.8489517, -2.2788111, -1.4320570, -0.5466233, -1.0093127, -2.8143455, 0.0880061, -1.3939994, -2.1272340, -2.2521977, -2.7402290, 1.7849308, -0.4821532, -2.2672026, 0.6809509, 0.9136314, -1.2411203, 0.3078890, -1.2197932, -1.4599665, 1.0066186, 0.4806967, 0.8629633, 0.6835951, 2.7766787, -2.4398540, 1.1223276, 2.2653617, -2.9274408, 2.9510369, -1.2871427, -2.9333855, -0.6912251, 0.8299761, -2.2340868, -0.2820885, -0.2780735, 1.7117476, 2.3300731, 2.4384339, 1.8596212, 0.7560404, 0.4714131, 0.3937447, -2.9107043, 0.9225049, 2.5850496, 2.2084493, 0.0404196, -1.2979969, -2.7759104, -0.6650872, 2.9569385, 2.7660146, 0.2321635, -1.8958140, -0.6221724, 0.6173596, 0.5518870, 2.0561694, -2.5989096, -2.3394210, 0.7540208, 2.7456593, -1.5916357, -0.4189588, -2.2412323, 0.2114440, 2.8166686, 0.5363482, -0.1511810, -2.4960748, -0.1781459, -1.8789793, -2.3701448, 0.3277580, 1.4847001, -2.6230044, -2.7372224, 0.8454972, 2.3963465, -1.4094941, 1.6984210, -2.1517965, -2.5881533, 2.6900178, -1.9025294, 2.8416590, 0.3667018, 0.1125374, 1.2715662, 0.3774072, 0.6269900, -1.7595931, 1.4072382, -0.3517551, -1.0376286, -2.6887607, 2.6901279, 2.8328959, -0.5245502, -2.5779251, 2.5698377, 1.5158323, 2.0799670, 2.5900657, 1.5024951, 0.3901550, -2.1256159, 1.3475663, 0.2905446, -0.4618245, -0.2892222, -0.1318619, 1.8771960, 1.7319434, 1.0826538, 2.5105219, 0.2593930, 0.8837335, 2.1544682, 2.4310635, -1.9684324, -0.4084282, -0.0790138, -2.6147280, 2.4645238, 2.1297089, -1.1730823, 0.9978720, 1.3609244, 0.7723116, 2.9903758, -0.9286971, 1.3896489, -0.2224370, 2.1883886, -0.4561498, 2.4722672, -1.3337490, -1.2880916, 2.9698236, 0.3234024, 1.3165134, 0.7820316, -2.3235964, 1.7587840, -1.0282488, 0.8225112, 2.4247555, -1.3009883, 0.0677655, -1.4512306, -0.2309304, -0.0501283, -2.1696346, -0.4150974, -1.5318028, -0.8888523, -1.4700186, -2.9824984, -2.9832381, 2.5909827, 0.8342039, -0.3499649, -1.1854091, -2.1794353, 2.9353661, -2.5817975, -2.4030629, -0.1208504, -1.3684464, -0.4948925, -1.3034197, 1.4834197, -2.9126643, -1.3590811, -1.2995521, -0.2871167, 2.7028470, 2.4000626, 2.3545412, -2.4955506, 2.9964422, 1.5913797, -0.8365839, -2.0766784, 0.6005996, 2.9830036, -1.4397704, 2.4209020, 0.0248218, -0.9063220, -0.7224452, 2.5861293, -0.2706737, 1.8732507, 0.6122651, -2.7524844, -0.1115900, -0.4553805, 0.1433230, 2.1318420, -0.5173890, 0.4631267, 1.0473971, 1.9043407, -1.0276248, 2.8222125, -2.9522655, 0.6704363, -0.6429993, -2.5538520, 0.7980070, 1.6137542, 2.2327877, 1.0232872, -1.6940046, -0.7709887, -2.6399282, -2.7212823, -1.0525675, -0.9852851, -1.2978458, 0.5811571, 0.6220806, -1.8238794, -1.6637259, 1.9953721, 2.2623720, 0.1883218, 1.8225440, 0.9305708, 0.1545184, -2.2743305, 1.7878328, -1.1642856, -2.4455324, 0.0687138, -0.9045417, 0.6490492, 1.0931038, 0.7326062, -1.8471137, -2.2396549, -2.1241951, -2.1594172, 2.7101524, -2.4020060, 0.1046685, -0.2548619, -2.8578138, 0.8284133, 1.7273646, -1.2231067, -0.3395657, 1.4333918, 1.1793799, -0.5263200, 0.9935715, -1.1185183, -0.6292723, 0.7955897, 2.9336269, 2.4728783, 0.1975981, 0.8331660, -0.7957811, 0.2812134, -2.5569996, -1.4959473, 2.8493068, -0.4801895, -0.4550216, 2.3462837, -0.1824604, 2.2513657, -1.7161377, -2.0035509, -1.8809259, -0.1415808, 1.3964937, -2.6106786, 0.3007183, -2.0964875, -1.6484838, 2.1207521, -0.2941439, 2.9942988, -1.9200118, -2.4077607, -2.9603830, 2.8226062, -0.4945194, -0.4075391, 1.3132249, -2.0846993, 1.4632744, -2.7474074, 2.1383165, 2.5771212, 1.8438199, -0.3867212, -1.5906492, -1.0511462, -2.0998910, 2.0792334, 0.8985657, -1.3760140, 2.0163631, -0.7747750, -2.3804056, 1.7506471, -1.1453419, -1.9296595, 1.3933301, -0.5732871, -1.8930773, 2.9268855, -2.4693500, -2.9015504, 1.0335266, -0.9336931, -0.5075208, 2.5646505, 1.9070730, -0.9414686, 0.2919791, 0.2623622, 1.9733510, 2.6029054, -2.4040627, -2.4022289, -2.6756673, -2.6513702, -2.2633634, 2.9289493, 0.9858347, 2.5069891, 0.1223218, -2.7312119, 0.5729070, 0.2227501, -1.7240361, 2.5300526, 1.9431138, -1.6686422, 0.6433860, 2.7505747, 0.7084125, 2.1827052, 0.3556727, 1.8125697, 0.2333074, 0.3419011, -2.0609273, -0.6925945, -1.7298540, 1.2454307, -0.0453321, -0.7767350, -0.3766626, 2.7283495, -1.6541300, -1.3076133, -2.1973873, -1.8370337, 0.2115611, -0.7766436, 1.2763019, -2.4418732, 2.0378013, 2.2137256, 2.2387238, 2.9679400, -2.3705624, -2.0891530, 2.5327437, -1.5445442, 2.1069851, 2.6039800, -0.9352225, -1.7965311, 0.0604660, 0.0549757, 1.2717425, -1.9540415, -0.9101819, 1.4502869, -0.2553140, 1.4785710, -2.6973994, -1.9454066, -2.9841233, 0.2122230, 0.9492835, -2.8958562, 1.2638547, 0.7579142, 0.9684121, 1.5849148, -0.8907476, -0.1667876, 2.2231303, 1.3911499, 1.3602387, -1.2037859, -2.5499982, 0.9678504, -0.9166227, 1.3925459, -2.3307224, 1.7187986, 1.7652912, -0.4557332, -1.5118502, -0.4787348, 0.8316217, -1.7107882, 1.0589515, -0.4963795, -2.5619548, 0.4819943, 0.3395253, -0.2904563, 0.5219247, 2.2555890, 0.8600572, 1.9697337, 1.1615924, -1.1866183, -2.5445596, -1.8892192, -2.6908841, -1.9819972, 2.0808990, -0.5217687, -1.4357245, -0.8990344, 1.6681618, 0.5377290, -0.2579209, -1.3924826, 2.6476152, -1.4380092, 1.6466885, 1.8783654, -1.9703571, 1.2819729, -1.9068660, -1.0473188, -0.2064249, -0.9598049, 1.0285053, -1.0528625, -2.2395834, -2.5589680, 1.0166883, -1.1694166, -0.6071352, -0.3651430, -0.5468669, 2.7346796, -1.0280442, 2.4388601, -0.1724921, -2.1780558, -2.0805180, -2.9012295, -1.2456498, -2.6629988, -2.4168873, 1.2869337, 1.1473340, 2.1957912, -0.1123008, -0.2166243, 2.9735020, 2.3182415, -2.9463725, -0.3350971, 0.6791466, 2.9113575, -1.1873728, -0.7249064, -1.4373110, -2.5271882, -0.6349053, -2.8380840, 1.7339352, 2.5614094, -2.9160567, 1.1838622, 0.1196644, 1.5180094, -0.0969802, 2.1901126, -1.9261236, -1.2007137, -0.5678436, -1.0982001, 1.4866453, 1.3362862, 1.7985583, 2.0389441, -0.2813462, 0.9740135, -2.0894341, -0.8982694, -2.5017078, -1.0594413, 0.3242815, 2.4018437, 1.3961793, 0.5276411, 2.4526743, -1.8029705, -2.5557935, 0.1929722, 1.4366284, 2.5486939, 0.4435588, 1.5009688, -2.0716430, -0.2579458, 1.7306934, 1.1432722, -2.0911855, -0.5184573, 2.3752423, -0.2545649, 2.9171169, 1.1801235, 1.4552794, -1.0149631, -1.1328450, -0.5725001, -2.6670203, -1.3386334, -2.2549768, -1.0735617, -0.8679722, -0.3601339, 1.4831705, -1.0316756, -2.1776066, 2.0512298, -2.5644616, 1.5055022, 2.5185648, -0.3991138, 2.3990441, -1.0315915, 1.6413227, 0.8718875, 1.4382906, -1.0732723, -1.1024351, 2.2410016, -1.6423973, 2.2884606, -1.0764106, 1.2523009, -0.1462424, 0.8415751, 2.8999787, 1.2356124, -2.1914687, 1.8417300, -1.0217173, 1.6857656, 1.1754480, 2.3881121, 1.5570773, 1.6817957, 1.9570736, 1.2770144, 2.3820645, -2.4740283, -1.3705813, 1.6669649, -0.0309142, -0.3347958, 2.2444165, -0.9782708, 2.5501161, -2.3537538, 1.2273385, 2.5260828, 1.9828311, -1.6367178, -2.1819798, 1.8458730, -1.0253994, -2.8348187, -0.2629145, -1.3879788, -0.6858342, -2.2140219, -0.3913233, -1.1657123, -2.4973702, 1.7701642, -2.4114297, -2.8754969, 1.4344196, -2.6022567, -2.9634197, 1.2036955, -2.8256044, -2.3967061, -0.6055660, -0.0514679, 0.3017889, 2.6175220, 0.2221549, 0.2141418, -1.2930370, 1.7821543, -0.2604659, -1.3918091, -0.4030735, 0.9021409, 1.8768485, 1.2776392, 1.5169066, 0.5900323, 2.2184152, -2.3058846, -0.8581945, -1.8326701, -1.3391321, -2.2964892, -0.7610347, 0.3470119, -2.1122304, -2.7265084, 2.5789441, 2.5445830, 2.1081519, 1.7477474, 2.6540146, 0.7170618, 2.0464928, 1.7295332, 2.1513669, -1.0208807, -1.1539701, -2.6501249, 2.2457523, 1.4892367, 1.7931516, 0.3920831, 0.8842752, -2.8803839, 2.1214892, 1.4269979, 0.7610666, -0.9365940, 2.6896983, -0.0005149, 1.9871832, -1.0565559, 1.9106242, -1.7102832, -2.1040451, -1.8849235, -1.0999348, -2.4347206, 1.4757279, 0.0308551, -2.8650175, 1.5424758, 0.4045877, -2.9313188, 0.3904400, 2.2487247, 0.5863210, -1.7371531, -1.7151631, -0.0665155, -0.0819494, -0.4940022, 0.1745180, 1.2625108, 0.8260612, 2.9109605, 1.1136985, 1.3326759, 1.5575267, 0.1855089, 0.8057686, 1.4063050, 2.4396089, -1.0929852, -1.2370765, 0.8923813, 2.0683964, 2.4315238, -0.8457471, 1.6684596, -2.2907132, -0.3858271, 0.3313162, 2.1439523, -0.2592952, -1.4536758, -1.2478835, -0.8261593, 0.2701783, -1.4275592, -1.6661872, 1.4057923, 2.5136967, -1.8560804, 2.2775025, -2.0408521, 1.8123595, -2.0245229, 2.1082446, -2.5869730, -0.0432532, -0.6681695, -0.9943764, -0.2781109, 1.6652938, -0.3159215, 1.0183114, 0.1271872, -2.4314844, 2.5327343, -0.1791725, -1.2952678, -1.9327397, -0.8510132, -1.0362470, 0.9385443, -2.8358021, -1.0017502, -1.2396051, -2.9598930, -0.4785821, -1.0806679, 0.6945293, -0.4073175, 2.8090320, 0.6385574, 2.0524281, 0.3844830, -2.3784946, -0.0253011, -2.1866026, 0.1511552, 0.1043418, -2.1621220, 2.2801775, -1.7086478, 2.7944305, 1.4690475, -2.2554940, 0.1509471, 0.3715651, -0.7154495, -2.5674861, 0.1879346, -1.5035890, -0.8597716, 1.0360380, -1.6586207, 0.1298420, 2.4506240, 0.4988685, 2.9670314, 2.5860903, -2.3515869, 0.1129031, 2.8133470, 2.6453901, -0.8944025, -2.2739167, -0.8193216, 1.2622149, 1.3725750, 2.9796490, 2.2151703, 2.2840062, 2.5828566, -2.6078659, 0.8202314, -0.3731492, -2.8439822, 2.8327858, -2.0670777, 1.0076398, -2.7795505, -1.4591098, 2.6435781, -1.2877473, 1.5686369, -1.1316031, -0.1903803, 2.1544071, -2.6852173, 2.0103724, 0.5320452, -1.7548924, -1.4891483, 1.3367313, -0.9609956, -0.9632301, -0.3147899, 1.1115299, -0.5611183, 2.6277178, 0.9253758, -0.8482254, 2.5311091, 1.7776811, -2.4652364, -2.1245420, -0.9047889, -2.7426410, 2.8195417, -1.5221989, -0.1832376, 1.6146291, -2.7165048, 0.3375367, -1.0013722, -1.5232293, 2.2866095, 1.1775613, -0.7716053, -2.0753522, 1.2918614, -2.8623299, 2.6872011, 2.3593330, -2.2977254, -0.5022952, -2.1614905, -1.4277151, -2.6434893, -1.1201664, 1.0187507, 1.6460404, 0.5402298, -2.2329665, -2.3428373, 1.4583674, 2.9906218, -2.7287336, -0.1121445, -0.9447654, 1.5458058, -2.7794480, 1.9386683, 2.8405828, -1.9968670, 0.2147492, 1.9175277, -2.0434695, -1.0975899, -2.3290019, -2.9024283, 1.1344701, 0.6125390, -2.4651458, -0.0185798, -0.0729588, -1.9994864, -0.3616760, 1.3774328, 2.4055171, 2.2335646, 1.6817208, -2.0020137, 2.3143376, 2.3155047, 1.8532417, -1.0155735, 0.5727665, -1.4639985, 0.2650831, -0.2038233, 0.7147274, -0.2022577, -2.8282933, -0.6562078, -2.6687814, -2.1823879, -1.0098703, 1.0782373, 2.2262110, 1.8103838, 2.5730857, 1.3428116, -2.6904327, 0.8720326, -0.1228412, 1.1834932, 0.1715367, -1.9939191, -0.8664241, 2.1935953, -0.0448417, 0.0395967, -2.4545179, 0.3095970, -1.2064633, 1.5121267, -2.2510568, -2.5893639, -1.9377232, -1.3389313, -2.0755499, -0.7794757, -0.5918331, -0.9915440, 2.9111198, 0.0310804, 0.1946558, -1.3020577, -1.3297026, 0.1837688, 0.3630524, -2.4177179, -2.5151327, -2.2981572, 2.1605658, -1.3139785, -2.5685054, 0.8684854, 2.6561083, -2.9776022, 0.7808754, 0.5442321, -0.3512144, -0.3711823, -1.5932116, -0.4865772, 1.9654117, 2.3706100, 1.8584626, 2.9340043, 2.0646393, 0.1834130, -1.0927139, 0.2205195, 1.1056937, -0.1192472, -2.4949100, -2.6402852, -2.6655671, -0.9930162, -1.3559632, 0.8642110, 2.3627742, 1.4638701, 0.3729091, -2.8555799, -0.3430501, 1.1955702, 1.6698634, 1.5568269, -0.1464866, -2.1947923, -2.2559088, -2.3358099, -2.0584439, -1.3724226, -1.6812519, 0.5324392, -1.1818109, -0.9504880, 2.9376776, 0.5143055, 0.6510152, 2.6966970, -2.1375322, 0.4115277, 2.5718912, -0.2344179, -2.6470454, 2.5505268, 2.7253957, -0.9548950, 1.6998271, -2.1505983, -0.8499747, -1.4362937, 0.5773782, -1.4218883, 2.8739241, -2.1754346, 0.1847934, -2.5543219, -0.2127801, -0.2658654, -0.5356166, 1.1511842, -1.3815561, -1.0052740, 2.1172287, -0.4856662, 2.9770931, 1.1252870, -2.7272123, -2.2467945, 2.4012475, -1.3832908, -2.0823033, -0.4928491, -1.8463683, 0.7925790, -1.6146586, -2.6973573, 0.6319514, 2.0688321, -2.0669568, 2.8245845, -2.7141731, 1.8425643, 1.8131700, -2.1476057, 2.1312738, -2.1000969, 2.6019037, 0.2986766, -1.9652618, 1.4760556, -1.3183097, 2.4903570, 1.0075730, -1.3278476, 1.1358299, 1.9044787, -0.4935857, 2.0736381, -1.5559718, -2.9198015, 2.5770851, 2.1170907, -2.1064626, 1.1321864, 0.9307310, -0.9108833, 2.6262519, -2.9554478, -1.4519278, -0.2768778, -0.8717010, 2.6198223, -2.9324185, 2.0832553, -1.6102553, -0.8198524, -0.9942916, 2.9247096, 2.8025751, -1.6751385, -2.6747444, 1.3155138, -2.3649202, -2.6922052, 1.0954308, -0.8784204, 0.8184565, -1.9974939, -1.9817760, -1.0221777, -2.8421481, 0.3535421, -2.2895219, 2.1615778, -0.8229014, 2.6192161, 1.5387701, -2.6416120, 2.8881165, -1.4882765, -2.9244348, -2.4346357, -2.5567324, 2.7734140, 2.8231373, 0.5419173, 1.7367899, -0.6265506, -1.1567864, -0.5578958, 0.6086312, 2.4267186, 1.5045457, -0.5810812, 2.8084296, 1.3880872, 0.0629018, 1.3995390, -0.7488571, 0.3340087, -0.1507612, -2.9435138, 2.1950902, -2.4552993, 0.9373229, -1.4898798, -1.5790818, 1.7574953, -1.6921555, -2.9734434, 0.7310881, -1.9278026, 1.0398751, -2.3781228, -0.3017756, 0.1081355, -1.6441809, -2.5225388, 0.7250142, 0.2035724, 1.4487655, -0.7340721, 2.1311824, -2.8427533, 0.2753081, 1.2032784, 1.5662001, 2.7744865, -1.1523525, -1.2718158, -2.2975698, -2.7666465, 1.2443467, -2.5778421, 1.7791558, -2.3157428, 1.0009140, -0.8810277, -1.9380984, -0.0088735, -1.6603645, -1.3852086, -0.7444181, -1.4209503, 0.0431379, -2.8723236, -1.0602541, 0.7606760, 2.1283753, -1.8375431, -1.6289643, 1.0783500, 2.1954701, -2.3770073, 1.5220025, 0.0506784, 1.2217113, 2.5917364, -1.6376278, -1.3661275, 0.1669888, -2.4886380, 0.8759607, 0.9461285, -1.9213086, 0.4633978, -0.1890766, 1.0660528, -2.6987495, 2.6742846, -0.6220754, 2.6170397, -1.4032178, 2.7056491, 2.2548009, -2.3516824, 1.3847708, -1.9974058, 2.3859059, -0.0573002, 0.2370180, 1.4678063, -1.7476929, 1.3051271, 0.7899720, 2.6487212, 1.3605510, 1.5268139, -2.5258597, -2.2976316, -0.5135043, 2.3678994, 2.5616868, -2.5553602, 2.0445047, 1.3838826, -0.3635730, -1.2536321, 0.6873258, 2.1252455, -2.0003866, 2.7573990, -2.0532917, 0.9350368, 0.4625580, -1.6788544, 1.0622865, -2.6143283, -0.2065245, 2.9147336, 1.6838553, 2.0099679, -0.9965663, -1.6002099, -1.1482677, 2.9496079, 0.1226484, -2.4957536, 1.1111219, 0.6428680, -2.7097243, -2.6508683, -2.5895075, -1.6289517, -1.8216745, 1.5260212, -2.9633047, -1.1173305, 1.4368823, 2.1987893, 2.1995206, 2.7127705, 2.4930514, -0.2223848, -2.6738035, 2.4046372, 0.2418986, 0.8830193, 2.3503718, 2.5581623, -2.1394688, -2.4193849, -1.7209090, 0.9553093, 0.7834867, -2.8229096, -0.1524026, 0.1086924, 1.5411561, -2.4461634, -2.2473406, -2.0565605, 2.2586428, 2.0300341, 1.6378823, -1.4659576, -2.8827429, 1.7637875, 1.2324202, -0.1483168, 2.7959591, -2.6176193, 1.4792854, -2.5757112, -1.7804207, 0.9595002, 2.4205276, 1.4343809, 0.0893154, 0.6928260, -0.7502546, 0.3771410, 0.6853259, 1.5832966, -1.4998329, -0.3320170, 2.2235219, -2.0347203, 1.2660158, -0.4801668, -2.6108148, 1.3848448, -0.7748491, 0.5756396, 1.9743384, 0.1935502, 1.8901028, -2.3291989, -2.6068043, 1.8100302, -0.2788941, 0.9413117, 0.7044195, 1.7809267, -1.3894111, -1.1840775, 2.4695663, 2.7801291, 2.3472749, 1.3262550, 2.4966746, 2.3032723, 2.5831713, -0.5742254, -0.6003725, -1.0066813, 1.2822442, 1.1642344, -2.7181989, -0.5622462, 0.7197465, 1.1466910, -0.1252596, 2.0867304, -2.0562003, 2.4206725, -0.7706040, -2.2623691, 2.3313173, -2.4370134, -1.9956048, -0.2205322, -1.5387735, -1.7337656, -1.8029513, 2.3567458, -0.8570442, -0.0694520, 0.7923130, 0.6625977, 2.2009450, 1.8048044, -1.7630706, -1.8364723, -2.7673741, -1.3214803, 1.2268574, -2.3226190, -0.5835496, -1.3464978, -2.5040864, -0.1161398, -2.1919214, -0.0954786, 1.2136809, 2.1831846, -2.5825742, 1.4429119, -0.3438570, 1.0954329, -0.3971498, -0.9290076, -0.0004401, -2.6729013, 2.9933254, -0.7412358, -1.9022367, 0.4667451, -2.3430557, 0.6400764, 2.5011044, -1.3894396, 2.9936903, 2.4222845, -1.8545327, 0.1804228, -1.7145517, 0.3531975, 1.5248648, 1.4417415, 0.8662420, -2.7911892, -0.7052132, -2.9802808, 2.8688510, 2.0833712, 2.1111077, -2.2929251, 0.0537109, 2.7932556, -1.6338919, -0.4035085, 1.9666174, -0.7051953, -2.4363929, -0.6922576, 2.1836884, -2.2572114, 2.8695630, -1.5795404, -2.8976604, -2.9151636, -1.2035382, 2.4989830, 1.5602429, -2.0173265, -0.5301660, -1.2498259, -1.2194401, 2.2558225, -1.6225529, -2.5201039, -2.1358202, -2.9660863, -0.5854276, 0.7703312, -0.5689928, 0.9307996, 1.3443786, 2.9321363, 2.9304572, 0.3758270, 1.9553885, 2.3830675, -2.9769355, 0.6022156, -1.1808142, -0.1926650, -1.8833923, 2.8196563, -1.1193686, -1.4566960, -2.5537502, 2.7619188, -2.0035655, -0.6843447, 1.1447637, -2.7544738, 0.4751631, -2.7455303, 1.8126797, 2.1044426, -0.4615311, -1.0167336, 2.4519544, 0.9599203, 2.4738544, -1.6806484, 1.3841778, -0.0614261, 2.6993948, -0.7254394, 1.0805557, -2.7358213, 1.1542277, -1.3203054, -1.8594958, 2.6200041, -1.2235783, -1.3259490, -1.7302053, -0.8903782, -1.3639324, -0.1059165, -1.9245965, -2.3584809, -2.2646049, -2.9790382, 0.8743968, 0.8130193, -1.8809434, -0.3816137, 0.4810576, -1.2218465, 2.3029330, -2.2105400, -2.1057567, -0.6633802, 1.2684882, -2.3033731, -2.7479027, -1.5665144, 1.7667240, -1.3019799, 0.8722906, 1.7402343, -2.1967285, -1.7316706, -2.2242260, 2.0708142, -2.0188622, 2.7781120, 0.7425466, -2.7059113, 2.9740509, -2.8747143, 2.1071984, 0.9619536, -1.5201199, 1.0979858, -2.2773656, 2.8572153, 1.0020032, -1.2557042, 1.6947604, -0.5376430, -0.4793314, 1.6088562, -2.4714893, -0.1606512, 1.8460705, 1.6594383, -1.2707165, -2.4111586, -2.0146687, -1.9756708, -0.7914095, -2.1570230, 2.2933313, 2.2735967, 2.6843559, 0.0285388, 2.6246228, -2.2147551, 2.6203617, -2.6100561, 1.1551546, -0.5641658, -0.8649631, 0.8256823, -2.8314617, -1.6859037, 0.7104420, 0.1326435, 0.3155531, -0.0178108, 1.0128806, -1.2084773, 0.7534649, -2.8648717, 2.2761346, -0.9952893, -0.1800060, 0.7874977, -1.6412891, 0.8038111, 0.4440473, 2.9154572, -0.9568380, -2.5802112, 0.0022756, -0.3065798, 2.9323778, 0.5876548, 0.4107791, -0.8136029, -0.2880429, -1.1260968, 0.8930379, 1.8279430, -2.0792069, 0.5435532, 2.8297452, 0.8846502, 0.4929997, 1.0379343, -0.8545677, -2.8262776, -0.6944988, -2.7972151, -0.9674180, -1.3076011, 0.4049720, -1.0613154, 2.7634399, -0.7065075, 0.7120147, 0.5849334, 2.2211445, -2.5238846, 1.1018930, -0.5746022, -0.3747537, 2.9793953, -0.4965329, -0.2904481, 0.9579050, 2.1165797, 1.0992451, 0.3604842, -2.4653301, 0.3071242, -0.1018337, 1.0549488, -2.6656628, -1.3625521, -0.4035355, -0.2406309, -0.5281896, -0.2740262, 0.9904101, 0.5826848, 2.8002443, -2.2541143, -0.4435269, 0.6561887, -1.1802464, 1.5707011, 2.5695524, -0.0825787, 1.5293742, 1.0367309, 2.7589934, -1.3549674, -2.9317446, -0.6902128, 2.5957169, -0.6758224, -0.1540176, 2.5449244, -0.8541402, -2.2997068, -2.3876435, -2.1362045, -2.5563359, 2.6524196, 1.3219368, -1.3127956, -1.3835349, 1.6590484, -2.6851736, 2.9407855, 0.5994417, 0.3140161, -2.4245489, -2.4354589, 0.9578557, -0.4806431, 1.1160066, 1.8113897, -2.0699889, -0.8757000, -0.2586717, -0.1180668, 1.6379425, 1.5462643, -2.5376318, 1.4258760, -1.9836884, 2.6896518, -1.4490629, 1.8933407, -1.1509055, -1.8423387, 1.2230107, 2.2695550, -0.0355880, -2.6393458, -0.4636108, -2.8779130, -0.3401292, -1.7128641, -0.4998840, 2.8813234, 2.2296482, 2.4672783, -2.2108711, -2.3924632, 1.8521902, 0.3753056, 0.6067515, -1.9593227, 2.8101761, -2.4662839, 2.3544294, 2.1431206, 1.7428576, -2.6167855, 2.2409223, -1.0939089, -1.3112040, 0.2612821, -0.0495499, 0.3015125, -1.9896460, -2.1597910, -0.1294893, 0.2358193, -1.5696546, 2.0312960, 0.3310815, -1.1960329, -1.1714168, -2.0585522, 2.7556397, -2.2741043, 2.7911868, 2.9449670, 0.2839936, -2.8314851, 0.4127898, -1.9244262, 2.5737911, -2.6252029, 2.8957746, -1.8378526, -2.9734496, -2.5555885, -0.6460400, 2.8749456, 1.0331255, -0.3129548, -2.3585503, -0.8386640, 0.9131838, -0.8428647, 1.1108806, -0.9072895, 0.9664911, 0.0695136, 0.2802003, -1.3518648, -2.8523288, -1.8574733, -1.1005880, 1.7615353, -0.9126384, -2.7594683, 2.1790980, -0.3207127, 0.0622847, 2.0602817, -2.4243789, -2.7022283, 1.4196881, -2.5329490, -0.0640924, 1.2933535, -2.6555841, -1.8040547, -1.5569630, -2.8353965, -0.2165941, 1.2250975, -1.5159069, 1.4878083, -2.8270198, 1.0176915, 0.4037889, -1.9890285, 0.7629358, 1.6014437, -2.5947624, -1.2091419, 1.3283207, -1.4579270, -0.7702169, 2.5988890, 0.4326838, -2.7674771, 1.3309370, -2.5951990, -1.0190344, -1.9515905, 1.5803105, 2.8600281, -1.6289595, 1.3134557, 1.3016531, 1.4475929, -2.3569976, 1.5461421, -1.0873571, -0.5849507, -0.1913396, -0.7990506, -2.7230821, -1.6190247, -2.0427483, 0.3502322, 2.0113144, 2.6582306, -0.4402904, 1.6801491, -1.2734241, 0.6399354, 0.9292038, -2.7453000, -2.9502868, -0.7906957, 1.6149908, -2.5053152, -1.2672284, -2.5085530, 2.7489850, 1.4178499, -2.3205720, 1.5587618, 2.7780576, -1.1853686, -1.4585208, 1.7857965, -1.7507807, -1.2754916, 1.6046464, 2.6967872, 1.8296284, -1.1638527, -0.2117775, 0.1975270, 2.9563513, 0.1336829, -1.5598214, 0.4783207, -1.5243288, 1.1238358, -0.2829117, 2.2290159, -0.8458393, 2.0479398, -1.6870136, -0.2091118, -1.5756549, -0.6929372, -0.8714609, 1.3772723, 0.0410375, -2.1918815, 2.4963094, -1.1465656, -0.5605821, -1.8790893, 1.4812357, -2.8473039, 2.0506348, 2.8937983, 2.0629017, 0.0566984, -0.6217841, 2.8826342, -2.1691537, 0.6634368, 2.7472937, -2.6300315, -0.0861840, 1.7440061, -2.4931875, -1.2677597, 0.8791176, 2.2785726, -0.6358975, -1.1057609, 1.0654451, 1.8375697, 1.9210281, -2.1213760, 0.4265947, 2.6785873, -2.2028196, 2.6380918, -2.2691158, -2.8696914, 1.5533579, 2.1792227, -0.0907158, 2.5933863, -0.7112965, 2.3656431, 0.7351160, -2.1161441, -1.1968609, 0.8114997, 0.8561967, 2.1530822, 2.9259301, 1.1079846, 1.1566809, -2.8220272, -1.1006329, -2.0044776, 2.4520641, 0.7320540, -1.4449997, -0.4910793, 1.4993461, 1.9704723, -1.1802937, 2.2965117, -2.3715351, -1.4420646, 0.9331719, -0.6970996, -1.0739767, 2.4501188, 1.4267987, 0.4368127, 2.4988659, 2.5449702, 2.6957564, 1.7237970, -2.0524658, -2.2424811, -2.7190370, 1.4018700, 1.6100265, 0.7433393, 0.5385926, 1.3460715, 2.9499784, -1.4972331, 2.8775791, 2.6801571, 0.1115962, -0.5076553, 2.8445700, -0.3547110, -2.4355628, 2.8085711, -0.1956734, -0.7099294, 0.0054092, 1.1513244, -1.8783442, -0.4698336, -1.4206978, -0.4086412, 2.9038295, 0.7296739, 2.2820329, -1.4650259, -1.4364986, 0.1703336, 1.8745227, -0.1487233, 2.3620342, -2.9838556, -1.2374903, -1.2121074, 2.1999460, -2.2700115, 1.6024116, -0.1423612, 1.1125841, -1.4188077, 2.9520158, 2.0236242, 0.4068511, -2.4470633, -0.9183608, -2.5340614, 1.2153299, 1.8200529, 1.5196373, -2.6218218, 1.2049105, 1.8579119, -1.7717958, -0.0495920, -2.7916898, 1.7968482, -1.3340484, -1.1352604, -2.7577748, 0.6039388, -0.9231145, -2.6503557, -2.7417924, -1.3502262, 1.3438776, 0.4415537, -1.4167920, -0.2109954, 2.0878339, 2.5210141, 2.2805064, -2.9293885, -2.4517725, -2.7495981, 2.6108560, -0.8911009, 1.4934127, 2.6517811, 2.1448908, -1.1373918, -1.4453850, -2.1466831, 1.0000347, -2.0253908, 2.7672998, 1.6189655, 2.9936835, -0.2599047, -2.7002549, 1.3337997, 2.5026414, -0.2638626, 0.3514005, -1.2541872, 2.5765479, 2.5155628, 0.5484489, -2.1312568, -1.9632954, 1.6608988, 0.7928360, -2.3575094, 0.1645589, -1.2716934, 2.5424478, 1.0368230, -1.1544762, -1.1298753, -2.8375798, -0.9441911, -2.2268195, 2.2033596, -1.9631706, -1.3935064, 2.3175273, 1.9209781, -1.8167061, 0.4654744, 0.9249996, 1.7857583, 1.0066608, -0.4754827, 2.5951132, 1.5268654, 0.8522096, -1.5848838, -1.6769679, -1.6223866, 0.9898638, 2.2421849, -2.5715047, 2.6902280, 0.8847069, 0.2954713, 1.2872965, -1.4281509, 1.4508283, -1.9506177, -1.3422480, 1.6773805, 0.6349926, -0.8261332, -1.1921923, -2.2300900, -1.3871091, 0.9824560, -1.9505106, 1.8112539, -2.4656271, -0.3677979, 2.6299302, -1.9771043, -2.3579753, -2.3015824, -0.6487862, -0.3260583, 2.9370812, -0.3796688, 2.0877592, -2.5556400, 1.9578133, -2.6315357, -1.8421238, 0.8412096, -1.3823799, 0.7774256, -0.6677448, 2.6883282, 0.5609620, -1.4668802, 1.1435038, 2.5676136, 0.9333331, -2.1824481, 2.9421522, -1.3159434, 1.1096597, -2.4308568, 2.9362213, 2.3005294, 2.9112523, -0.5548237, 2.4736760, 0.8234591, -1.7576428, 0.2311943, 1.5293473, -0.2718800, -0.9902330, -0.2675725, 0.1912849, -0.1000799, -1.4359984, 2.3770191, 0.0971124, 1.0902430, 1.1441258, 0.3285317, 0.2110269, -1.6698519, 1.3492236, 2.3332027, -0.6093328, 0.9763373, -0.3787144, -2.0910803, -2.0009857, -0.4999366, 1.3254934, 1.2954296, -0.3909579, 1.1954102, -2.0925670, 0.5908926, -2.8144450, -1.3767406, -0.2277149, 1.6475723, 2.3310949, -0.5051299, 2.1165637, -0.0456829, -2.9018001, -2.8480404, 1.5186237, -2.6912983, -0.6782256, 0.2000163, -0.2259045, 0.3406461, 1.8700968, -0.8000331, 1.7058305, 0.6551541, 2.2563618, -2.6614001, -1.4971251, -1.8574491, -1.0747857, -1.7873875, 0.1402519, 2.6421187, 1.2190694, -0.0296710, -2.9626540, 1.4097833, 2.9736999, -1.4226468, -1.2616040, -1.6041606, -1.7802425, 2.2791849, 2.6141836, -1.0258761, 2.8629898, -2.0205115, -0.6710059, -2.6620654, -2.1897397, 0.3030567, 0.1547266, 1.7786772, 2.9988962, -1.6890003, 2.0333459, 2.8293393, 1.4729968, 0.2773837, 2.4905652, 1.0492949, -0.9573837, -2.1897974, -2.2887543, -0.2438752, 0.6126073, -2.6241130, 1.2423803, -2.0618430, 2.8160534, -0.1833627, -0.2761407, -0.2607385, -2.9229096, 1.8143413, 0.9920238, -0.1895342, 0.2496843, 0.4156337, -0.4129266, 1.4981899, -0.0833091, -2.6867030, -0.9197416, 2.0464538, 1.9288691, -0.3009736, 1.9258509, -0.8180040, -2.5387040, 0.2470880, 2.5744869, -2.5186522, 1.6684624, 1.8223773, 1.5643095, -1.5414828, -1.2201202, 0.1856749, 2.2621380, 0.5830643, -1.2343409, 0.6530387, 2.0941427, -2.4325511, 2.4948864, 0.6672031, 0.9207761, -2.9083260, -1.0809526, 2.1425663, -0.6354450, -2.6031468, 2.5365744, -2.0928219, 1.8429422, -2.5739911, -0.0991637, 1.2340546, 1.8959960, -1.9043059, -0.6693825, 1.2415684, 0.2598134, 1.1636811, -0.7740796, -1.5603310, 0.7852282, -2.5541335, -1.1241552, 0.0440543, 1.1982941, -0.3879077, -0.3036915, 1.6041354, 0.1529127, -1.7627537, 2.1228159, 0.2946977, 1.5501126, -0.1292458, -2.3571567, 2.6863231, -1.6344466, 2.4749644, 1.9178296, 0.3048203, 1.3321111, 1.2558117, -0.2752455, -2.3292181, -1.0717395, -2.2158820, 1.3675387, -1.3980824, -2.3221360, -2.0619038, 1.6641686, 1.7989319, -2.2375746, -0.0807435, -1.1890748, 2.9268463, 2.2593321, 2.1737336, 1.6420025, 1.9588063, -2.4059407, -0.9067161, -2.5814596, 2.2289676, 0.3238035, 2.8320071, 1.8220390, 2.8375128, 0.9177905, 0.0074081, 1.4748021, -1.4490418, 2.6100973, -2.7281737, 1.2999543, 0.4063791, -1.2481273, 1.0551817, 1.3510216, -1.5002528, -1.2187796, 0.9864547, 1.1271361, 2.0235571, -0.6526821, -2.1118778, -1.2353758, -0.9615100, -1.9114336, 0.2302034, -1.0307007, -2.2421915, -2.1524881, -1.5635283, 1.3240677, 1.0305389, -1.0991601, 1.5226755, 2.6007261, 1.0137534, 2.2168331, -1.2243320, -1.7333985, 2.3189009, 0.1781770, 0.8367562, -1.9593571, 0.3625807, -2.4000654, -1.8086000, -1.3401662, 1.4243435, -1.7064166, 0.0398081, -0.2193919, -2.3444918, 1.3200174, 0.4363449, 2.9952413, -2.3973390, 1.9864608, 0.6129185, 1.6121146, 2.4997873, -0.8911528, -1.1638473, -0.8783993, -0.1758937, 0.9861215, -0.1313288, 1.4344808, 0.5031243, -2.6611464, 1.2501905, -0.5505617, -2.0704859, -2.5726237, 2.9398256, -2.7799268, -0.9722779, 0.0479190, 2.3599845, 0.6659583, 0.3623674, -2.3561440, -2.7531413, -2.0473790, 1.6896588, 2.3769579, -1.6300849, -1.1408073, -2.9976142, 1.8068621, -2.0900524, 2.2773524, 1.3948748, -1.6756576, -1.0533463, -0.5609333, 2.1576474, -1.9848267, -1.9953383, -0.1229028, 0.1175117, -1.0296671, 0.7394158, -2.5135836, 1.2826213, -1.4261629, 1.5439779, -2.8475178, 1.1097474, -2.0432367, 0.2566169, -2.8938244, -0.1325770, 2.4187124, 2.1829898, -2.4235228, 0.3488555, -1.9758360, -2.5060300, -2.9156038, -0.6083634, -2.5539220, 1.9104516, -2.4574712, 2.9460915, -0.5120889, 2.3294075, -2.2266770, -1.6041071, 2.3534440, 0.1699672, 0.5439340, -2.4573293, 1.3588076, 0.1009578, -1.2108662, -2.8214559, 0.0459369, 0.6536504, 0.1791752, -1.7667264, 0.9475103, 1.1998030, -2.9579476, 1.1381043, 0.9561582, 1.5799673, 0.7394445, -0.2853649, 0.7655699, -1.0136106, -1.8492896, -2.0169160, -0.9865032, 2.1477261, 0.6861279, 2.0263584, 2.3579175, 2.5095631, 1.4324435, -2.0203656, -0.8230641, -1.2682069, 2.5931383, 2.5884065, -0.4217536, -2.9315098, 1.1285907, -0.1967494, 1.4349836, 1.2059397, -0.7438644, 1.0837430, -2.1373603, -1.5837610, -0.8979739, -0.9549511, -2.0135205, 0.1472058, -0.7281174, 1.9588397, -2.7135157, -2.9369795, 2.6657070, 0.9973213, -0.9598558, 1.3526444, 1.2694047, 2.5673053, -0.8254513, -1.5786756, 2.6647682, -0.6742181, 0.8334949, -1.3499200, -0.9372361, -0.4231000, 2.4556017, -1.3761272, -0.6292117, 1.4950582, 0.0735591, 2.9749329, 0.7221066, -2.7176513, -1.8838295, 2.3660293, 0.9905572, -0.9842869, 2.7224177, -0.7495854, -0.8509975, -1.9141955, -2.0466332, 0.9676488, 0.8008467, -1.4483420, -1.4894787, -0.5204098, -1.6055392, -2.5701524, -0.7714275, 2.1670216, 2.4599502, -0.0548801, 0.9783733, -2.9972429, 2.1953003, 2.8374195, 2.7346287, 2.0027317, 1.8795145, 2.4149689, 1.1963310, -1.4285310, -1.7279550, 2.2033686, -0.8023272, -0.9330612, -0.5093010, 2.9829112, 2.5152277, -0.7094183, -2.6115759, 0.8818772, -1.2136437, 1.4482258, -0.2007853, 0.3492919, -1.4961613, 0.3993254, 1.1872107, -2.5245067, -0.5899087, 2.2248276, 2.7166686, -2.7015096, 2.9520459, 0.3030075, -1.4741430, 0.6868371, -2.9576446, -0.4003389, 2.8412626, -1.5392235, 1.0241778, 2.6600604, 2.6831991, 0.1894700, -0.2381333, -2.2866471, -2.7312081, 2.6780474, -0.5914083, 0.8941353, -0.7575674, 1.9736024, -1.4424730, -0.0475658, 2.9348019, 1.6979960, -1.4581239, 2.6182310, -1.4284925, -0.6662386, -1.9384453, -2.1404986, -1.5805884, 0.7047830, -2.5334295, 0.6060339, -2.7845602, -0.6613408, -2.1742448, -2.9746791, 1.8167462, 2.4334973, 0.3359029, -1.8289296, 2.6789012, 0.2259312, 0.3548455, 1.1655642, -1.7071519, -0.3687508, -1.5878730, 0.8485586, -2.0856791, -2.7331013, -1.7669559, 0.3975381, -1.2242071, 2.5742808, -2.2356316, -1.6130414, 2.0118173, -1.9611746, 1.3482893, 0.2320292, -0.9699043, 1.0158583, 1.7643098, 0.6731198, 2.5293898, 2.8762647, -1.0552524, -1.1377023, -2.7538456, 1.5564798, -0.7964809, 0.0790590, -2.9934511, -1.9197749, -0.6661771, -0.3673835, -1.2184774, -1.4962750, 0.4893598, 2.3376529, 2.0899884, 0.5812831, 2.5447502, 1.2504410, -0.7809342, 1.8118779, 0.8749400, -0.6475259, -2.0994452, 2.9246689, 0.5586559, -0.8007405, -2.1908851, 1.2040484, 1.7166485, -2.3975199, -0.0581689, -0.1464031, -0.2395373, -1.0446429, -0.7027466, -0.1142316, 0.1359510, 1.8048472, 0.8727554, -2.1295737, -0.0856964, 1.1502358, 0.2379057, 1.1787422, 0.9480273, -1.6479932, -2.5227294, 0.1302975, 2.4301383, 1.4248009, 2.7953023, -0.9443029, 1.0630909, 2.7516201, -2.6516178, -2.2838851, -0.1384185, 2.7472304, 2.7440633, -2.3716336, -0.9862099, 2.0538719, 1.6174886, -1.6308601, 2.8696444, -2.1057737, 1.6172009, -2.6918593, 1.3187796, -0.0929262, 0.9538396, -0.1009516, 0.6681969, -0.2082916, -0.6426009, -1.8552293, 2.5415264, -2.2274939, 2.9077998, 1.6265715, 1.2930745, 0.2119647, -0.8010443, -0.6235555, -1.3321031, -1.7564126, 0.0532910, -0.6853093, 2.4636395, -1.4133556, 1.9142605, -2.7101863, -0.7021834, -1.1842779, 1.6404260, 1.9919340, 2.9548066, 0.9237237, 1.8116234, 1.6007849, 1.2821383, -2.8656897, -0.0945105, -0.6042729, -2.3307616, -1.5174350, 2.4715262, -1.8687515, 2.5393819, -0.9285511, 2.1835282, -1.0154420, 2.7352495, -1.6060915, -2.4709496, -1.7100787, 1.3303337, 1.7511609, -2.0906664, -2.7193328, -1.2933614, -2.1458202, -0.5729738, -2.3788632, -0.8343251, -0.3259823, -1.3475140, 0.0807992, -2.7462409, 1.5096951, 1.1979192, -2.6202731, 2.7701923, 1.7552228, -1.0973692, 0.6897969, -0.5607567, 0.7555953, 0.0093942, 0.4179274, 1.7674947, 2.2038658, -1.4598518, -2.3861078, -0.6807673, -2.7109806, 1.4235419, -0.0522188, 1.2700675, -0.5944995, 1.9295292, 1.8012555, 0.6616642, 1.2527731, 0.6585718, 0.5656344, 2.4667011, -0.7943379, -1.0257187, -2.7407014, 2.0883909, -2.5622203, 0.6004658, 0.4839886, -0.5787179, -2.2988440, 1.0239979, 1.8738051, -0.7429908, 0.6431525, -2.0122339, 2.4090668, -0.1106574, -0.7961747, 1.8978453, 0.9254303, 1.7075298, -1.3097423, 2.3159687, -1.3868370, -1.8720229, -0.5174073, -0.0689688, 0.2742193, 1.8113139, 0.3176768, -1.2120350, 1.8478120, -0.4295878, 0.3634222, 1.8775778, 0.5933253, 1.9421321, -1.4109285, 1.7957541, 2.5012708, -0.0043927, -1.5030729, -2.5063561, -2.1925835, 0.8772890, 0.9689016, -2.2844982, 0.3790415, 0.1236368, 2.4891264, -1.1988471, -1.0652530, 0.6619812, 1.8976820, 0.5029040, 0.3558135, -1.6334840, -1.0724554, -2.2690827, 2.7889365, 1.2216077, 0.2554366, 2.8529330, -0.0686303, 0.6126789, 0.2230877, 2.6432581, 0.2994384, 1.4571215, 0.6684477, 2.4508887, 1.1469077, 0.6588594, 2.1924117, 1.9690514, 2.4214811, 0.9362738, 1.8281745, -1.2782718, -0.2131736, 1.7344236, -1.1022269, 2.9906092, -2.0173523, 1.9127721, 1.9872413, -0.2277402, -2.8815415, -0.2081868, 2.8908529, -2.5386740, -1.6364486, -2.2023760, -0.1401172, 0.5227815, 0.5873062, 2.6705271, 0.3708922, -2.8710910, 1.8462375, 0.1351162, -2.5618837, -0.9494132, 0.3883501, -1.9712944, -0.9586677, 1.7237954, -2.3502852, -0.6785800, 1.8114787, -0.5995715, -1.9020835, 1.9612558, 2.1572003, 1.5839020, 0.5837522, 1.0299879, 1.0053060, 1.4140223, 1.4884214, -2.3419761, -2.9856989, 2.0948104, -1.4432065, 2.7537443, 2.6976926, -0.4178034, -2.2507033, 2.1532051, -1.9061965, -1.6315653, -2.1222960, 0.7413045, -2.6991686, 2.7670669, -2.2364284, 2.9697222, -2.6464377, 1.9497347, -2.2246744, -1.4358503, -2.3619078, 1.3530055, -1.5468543, 1.1125587, 2.3599185, 0.6201609, -1.2027822, -1.0649284, 2.0419711, 2.0670548, -1.0177923, -2.3845286, 2.6080334, 1.4817854, 2.9579395, -2.5615934, 1.2768138, -0.0290848, 2.7101434, -0.5876228, -1.1655153, 0.8392208, 1.2736468, 1.5132341, 2.9707125, -2.8576588, 0.8988487, -0.4871611, -0.7451406, 2.4137700, 2.1003856, -2.5684093, -0.5808836, -1.4531081, -0.5406771, -1.0791615, 1.2357899, -1.7585910, 1.0627419, -1.4394160, 1.7430533, -0.8346123, -2.5020216, -2.2573375, 0.4695721, 2.4545538, 2.5293221, 0.5619575, -1.5733870, 1.1772519, 0.3635764, -1.7030356, -0.7733475, 1.5521816, 2.3000584, -1.3946335, 0.8486229, 2.0717213, 1.4752375, -0.1030468, -0.3915947, 1.0274102, -2.2063255, 2.5384941, 2.4578085, 1.2025004, 2.4169866, -1.9692301, 0.2993863, 0.0463170, -1.8949436, 2.5298647, 1.7070882, 2.6863968, -0.7449014, 0.0135791, -1.9488813, 2.3249464, 1.7357998, -1.9205341, -0.5289005, -0.2363527, 1.8390760, -0.6683446, 0.5268482, 1.6522576, -1.6727396, 2.6949544, -0.2121289, -2.8154129, 2.9874768, 0.0405222, -2.3025800, 2.2696466, 2.2699318, 2.0009741, 2.9691033, 1.3558903, 2.6951284, 1.1053400, -0.6764215, 1.1031273, 2.8370958, 0.3372160, -2.3667717, 0.6293143, -1.4815613, 0.4167883, 1.1540179, 1.8852450, -0.1287819, 1.4853533, -0.9380841, -0.8816541, -2.9929377, -1.7989096, 2.0983506, 2.3538246, 2.6989572, -1.3448455, 0.5586830, 1.2447040, 2.0178523, -2.9637925, -0.7800807, 1.4648551, 1.5047184, 0.3019717, -2.6414784, -2.6662394, -0.5095949, 1.7694073, 1.4181313, 1.3228852, -0.9876803, -2.3421790, 0.3222284, -2.4813692, 0.0301586, 2.9973767, -1.3188420, -2.8931211, -2.7400006, 1.9727885, -1.0588229, 1.0130340, -0.4514502, -0.2843971, -1.7691901, -1.8769859, -1.8961061, 0.3724187, 1.5966436, -1.7928626, -0.9364250, -0.2001862, -2.8616818, 0.8857276, -2.9219856, 1.3996577, -2.5554310, 1.1549180, -1.3032069, 1.4336682, -1.7468045, 2.6359152, -2.1730373, -0.2092296, 0.2296345, 2.9471488, 0.3501169, 1.5699874, 2.0784537, -1.4543908, 0.0705399, 2.3111449, -0.4869171, 2.6109859, 1.3920305, -0.4030019, -0.3082508, -0.3922167, -0.6216964, 0.3750841, -1.0883669, 1.7482748, 2.7200293, 1.9280406, 0.4964557, -2.9375309, 0.3252373, -0.1097725, -0.8090665, 0.6216294, -0.2434173, 2.0475460, 2.8170401, 2.9364096, -0.6457290, -1.3861683, -2.7485196, 1.8929609, 1.6759162, 2.2710186, -1.5243893, -2.5704686, -2.9738278, -2.3034074, -2.0072942, 2.1415135, -0.0383746, 1.2581506, 1.4716634, 1.9003651, -1.9499062, 2.0491941, -1.3152481, -2.2394471, -1.2937501, -0.9670002, -1.9095824, 2.7503599, 2.9409161, 1.7429907, -1.6652089, 1.8425926, 1.5648882, 0.2018551, 2.4426510, -0.6789840, -1.7315660, 2.6947186, 1.1469594, 2.4086590, 2.7216842, -2.0902809, 0.8218999, -0.7781895, 1.0764980, -2.3056071, -1.0969431, -1.7410135, -2.2560995, 2.5239832, 0.8283234, 2.5900668, -1.8209906, -1.3847367, -0.8286398, -0.5813845, 0.0756613, -2.3926333, 1.3937508, -0.2200622, -0.6654671, 1.4798992, -1.9894435, -0.6343504, -1.7788143, 0.9010789, -1.3881078, -1.8676494, 1.5900613, -1.5354339, -0.5080747, -1.8979166, 1.1067348, 2.5313136, -1.9485949, 1.2088244, -2.4633699, 0.0683961, 2.5242405, 0.8060949, 1.2432047, 2.1982999, -0.3283216, 0.1968316, -2.7612973, 0.6812924, -0.2332562, 0.7712162, -0.5615220, -0.8245845, 1.5726441, 2.5057956, -2.6894156, -0.8763053, 0.9137804, 2.0902376, -1.4560561, 0.1533671, -1.3531986, -0.0973405, -1.5340300, -2.3806682, 0.2704262, 1.2808334, 1.1264338, -2.3834554, -0.4524227, 2.7738579, -0.4064429, 0.3404370, -1.6437232, -2.3769884, 2.4538428, -1.6203375, 0.5982439, 2.2377179, 2.9432414, 1.4422546, -0.9756417, -0.6321741, 2.7258139, -2.2314719, 2.6664619, -0.1311824, 2.6580039, 2.5085315, 2.7415741, 1.3701427, -1.0263521, -0.2638369, -0.3404236, 0.9172880, -1.3574959, -2.8849938, -1.4313321, 1.7353175, -2.1416292, -2.3635519, -1.4372756, -1.5349697, -0.1191404, -1.7251180, 0.1648209, -0.8166581, -0.8080226, -0.6210463, 0.1719246, 2.6070419, 0.7500825, -2.4033105, -2.3242606, -0.3387124, -1.6443281, 1.1261741, 1.0224332, 2.5896899, 1.7247672, -0.8152708, -0.4726073, 0.8597564, 2.4522407, -1.2293560, 0.6747918, -1.1870577, 0.7644721, -1.0910483, 0.9768590, -2.5367227, -0.9450981, 1.4999063, 1.0697955, 0.0927648, 2.3738435, -1.2433703, 2.8698964, 1.3831577, -0.9821302, -1.9249697, -2.9673170, -2.0431243, -0.9062035, -2.9393386, 2.2709824, 1.6770810, 1.7109299, -0.4015096, -1.4119578, 2.8364297, -0.0976709, -0.8524891, -2.1128856, -1.2767434, -0.1501717, 0.7471072, 1.7623011, -1.5160275, 2.5796571, 0.0737259, -2.9921622, -1.4381092, -0.2809915, 2.6370888, 0.1918868, 2.1927787, 0.5805763, -1.0035718, 2.1057837, 0.2229337, 1.8743675, -1.9101212, 2.7193744, -2.7646375, 2.5915353, -1.1271703, 2.6168322, 2.9819510, 1.9166445, 0.7689786, 1.7453635, 0.3112899, 1.7680362, 1.1438616, -1.9668779, 0.7984577, 0.6976562, 2.7223067, 0.8756045, 2.2524546, -0.3163828, 2.9131991, 0.5921055, 2.5322724, -2.1612752, 2.8882967, -1.9088779, 1.4298753, -1.2724437, -2.6085470, -1.2902728, 2.2886971, -2.7731542, 1.3043192, -2.8497292, 2.8968513, -0.9671175, -0.6346372, 0.4094442, 0.4318263, 1.5642340, 2.8468648, 2.2373418, 2.5580600, 1.1084734, 0.4025870, 0.6353699, -0.2519483, 0.2604904, -2.3846319, 0.7380913, -1.4345515, -1.9199519, -0.1709221, 2.8006967, -0.2617183, 1.2815276, -1.1603607, -2.7666347, 2.5720184, 1.6980644, -0.5129700, -0.0701834, -2.2451478, -1.7636953, 0.4938137, 0.3730028, 1.6295326, -1.1912056, -0.1510105, -1.1430835, 2.4711390, -0.9251857, -1.3736723, -2.6976637, 2.3662108, -0.1426096, -0.0341544, -1.4452036, 1.1880735, 1.2842192, -1.9251913, 1.1456762, -2.7187493, -0.8017838, 1.5151977, -2.6136803, -0.5895505, 0.0463244, 1.4560336, -0.9544518, -1.5504779, -2.3123060, -2.5122417, 1.2364479, -1.3429908, -1.6070043, 1.0306417, 0.1560774, -1.5515494, 0.4908575, 1.1201915, 2.7228506, 1.3400742, 1.6972200, 0.0461776, -2.6301147, 2.3197876, 0.6385069, -2.3227438, -2.2549116, 1.8913713, -1.3921638, -2.3984105, 0.3705548, -1.5169554, 1.8356721, -0.2512835, 2.0081848, -1.7602646, 1.0329428, -1.4643050, 1.1877042, 1.6050719, 0.4548951, -1.9332555, 1.3450655, 1.5635048, 0.3461770, -1.4832588, -2.8557202, -1.3349879, 1.6504048, -1.2846764, 1.5792712, -0.2629427, -1.5441189, -0.5466113, 2.8551112, -2.1715001, -1.1946570, 2.1034967, -2.7636103, 2.9685041, -2.1308080, -2.5498313, -2.6419688, 1.1618646, -0.6995263, -1.4275378, 1.3930656, 0.9517999, 0.7341352, 2.5800041, -1.5893875, -2.0068362, -1.0186806, 0.5641496, -2.8637025, -2.1961193, 1.3796792, 0.5712655, -2.7480470, 2.6182951, -0.2016989, 2.7088118, 0.6890784, -0.6531870, -1.3166223, -2.4274197, -0.3940246, -0.2943527, -0.2612535, -1.7789659, 2.6342937, 1.2312166, 2.6234876, 0.3091881, -2.0886628, 0.3914723, 2.4619890, -1.4808292, -0.7801174, 2.2605669, 2.3789266, -0.1227129, -0.7086448, -2.1350361, 0.6072603, 2.2150753, 0.1641213, 0.1163389, 2.5954404, -0.5602774, -1.3367172, -1.7549858, 0.6048661, 2.3454575, 0.1014981, -0.5263914, -0.4540699, -2.8814349, -0.9456093, -2.4238502, 0.0903966, -0.3970383, 0.4780366, 0.9892551, 2.4641025, 2.1939260, -2.9705464, 1.5965823, -2.5552962, -2.5006457, -2.5440190, -2.2965685, -0.6948890, -1.9127247, -2.6991520, 0.0961099, 2.6899699, -1.3974685, 0.8099574, -0.4490807, 2.7214899, 0.7412240, -0.7925006, -1.2041097, 2.1476010, 2.1503126, -1.7589175, -1.7124729, 2.6359872, -0.2156731, 1.7586610, -2.3787651, 0.4346598, -1.8665552, 2.1120167, -0.6167547, -2.9662790, 1.4614183, -1.6926935, -2.4402178, 2.6987879, 2.2171526, -1.4335945, 0.2268906, -2.5809429, 0.0414328, 0.9149110, -1.8786649, 1.1991529, -2.5955279, -1.7465852, 2.8606461, 2.4733809, -2.5636483, 2.8086033, -1.8562573, -2.3000664, 0.8065845, -0.5507937, -1.2800531, 0.3182178, -1.4096672, -1.6633489, -2.0462657, -2.6806735, -2.4594449, -1.8212247, 1.0294605, -2.9742590, -0.8329707, 2.2262038, 2.9942108, 0.1511197, -0.0702830, -1.5948325, 1.3430199, 2.3954214, -1.9819242, 1.5714929, -2.5635828, 0.2466356, -0.3665978, 2.4219275, -0.7119192, 2.2068304, 0.6539402, -0.2120807, -2.1174634, 0.3096532, 1.6215913, 0.3375743, 1.0809442, -0.5440515, 2.8339321, -2.2861963, -0.5326844, 2.0296567, -2.1343291, -1.0682916, 0.6686787, 0.0479496, 1.5467411, 0.7575443, -2.8634740, 2.6136610, 2.0581912, 0.0320819, 2.3127826, 0.6696695, -0.9444699, -1.0801453, 1.4091367, -1.7573271, -0.8130138, -0.5684477, -1.7209559, 0.3699770, -1.8459547, -2.9144714, -2.8352398, 1.5909854, -1.8932330, -0.9283645, 2.4013069, -2.2556897, 1.7760920, 2.2675147, 1.0591899, -2.5776629, 0.6248420, -0.2813571, -1.2607683, -0.6554490, 2.4132482, -0.0914649, -1.1120556, 1.3456167, 0.1195136, 0.4462410, -2.3562386, -0.1707408, -1.0604702, -2.0000016, 1.2862063, -1.9875185, 1.0922857, -2.4819305, 1.9502219, 2.3923564, 1.3559986, -1.7012292, 2.0637841, -2.8544230, 1.8900048, 1.6739074, 2.3674648, -2.1118334, -1.1900195, -2.9493120, -1.7308301, 0.2825989, 2.7254854, -1.5912851, 0.0766466, -0.1699209, -0.3639688, -1.6090110, 2.8650145, -0.6302551, -2.5315141, -1.9311190, -2.9461263, 1.4879006, -2.2327750, 0.8905650, -2.2316648, 0.1832579, 2.7537129, 1.3084152, 1.9818057, 2.6571235, -2.3481290, -1.5397942, -1.6937670, 0.4478371, 1.3239260, -0.9561457, 1.7744843, 1.4184649, -1.5525357, -0.8027819, -1.2915361, 0.6229948, -0.1049604, 0.3936277, -0.7345639, -1.6235057, -0.0290470, -0.5666983, -0.0277354, 1.1879748, -1.4409820, 1.6250944, -1.4054719, 2.6707139, 0.4310584, 2.9063388, 1.5242768, 1.1703159, 1.5657007, -2.4429452, 0.6021541, 0.4772359, -0.7094894, -2.8262965, 2.4971734, -0.8765248, 1.8499561, 2.4166376, -1.2477994, 0.3690813, -1.0218246, 1.9478965, -2.5581263, -1.8737264, 1.6604631, -0.3760260, -1.0689602, 0.1759576, -1.2299608, -0.9240652, 0.4198546, -2.5215878, 0.9290924, -1.5154490, -2.2810018, -2.6065385, 2.8491403, -2.2534982, -0.5824086, -1.2624916, 1.5901764, -0.8404630, -1.7773371, 1.4242800, 1.1678187, -0.6888041, -2.2140665, -0.3715741, 1.9642653, -1.2829883, 1.5238361, -2.4583766, -2.1499436, 0.7176010, 2.2233436, -2.7451912, -1.7701290, -2.1210618, 2.6838912, 2.0307963, 2.2354570, -1.1166541, -0.5491637, 1.7475731, -2.6574923, 1.7435313, 1.3387916, 0.1009325, 1.1868332, -2.6431130, 2.1598057, -2.8054540, -0.7669262, -2.4285093, -1.1086380, -2.9542808, -2.9334213, -2.1228308, 1.3518485, 1.5886077, -2.7610631, 1.6162624, -1.5076050, 0.7072872, -1.0082920, -1.2081265, -1.3611938, 2.2014150, 0.6090918, -0.9276433, 0.2382676, -0.5294441, 1.3772594, 0.7808640, 0.8746281, -2.2855646, 0.7965599, -2.4567019, 0.6174570, -1.1883009, 0.8007935, 2.3205632, -0.2754342, -1.8446423, -0.4351971, 0.4998578, -2.6860932, -0.9434962, -2.8274650, -0.9359373, 2.6725117, 2.4276806, -1.3168285, -1.5894740, -1.3888388, 2.8711189, -1.2896563, 1.4126103, -2.3890558, -2.2555679, 2.1011428, 2.0436106, 0.4280769, 2.7861282, -1.7364916, 2.1192987, -0.2698652, 2.4988037, -2.8660555, -1.2696006, -0.5017769, 1.6679480, 0.9429256, 2.7878609, 1.8611986, -1.8515398, -2.7623074, 1.3029922, -2.8201589, -2.7306529, 2.7873743, -2.0598800, 0.3604035, 2.7294368, 0.3127539, -1.0444562, -2.4945070, -0.3069345, 0.2495654, 1.6677167, 1.8443119, 0.8819934, -1.0998485, -2.7083191, 0.5303112, -0.0241769, -0.5534860, 0.1581904, 0.3459676, 0.9104774, 0.7369970, -0.0144912, 1.5004369, 2.5857336, -1.0405018, 0.4790480, 1.7393392, -0.5049726, -0.1933041, -2.2582391, -2.9689514, 0.5072212, 1.6171378, 0.6599660, -2.7667899, -2.7451540, -1.4859553, 1.4267842, -2.9686176, -1.9445603, -2.1914353, -2.1704920, 0.7963844, 0.1383718, 1.9919760, 0.2580539, -2.3751782, -0.5744282, -0.7777295, 0.8985036, 2.2162683, 0.1717986, 1.0136916, -2.8531507, 2.5256595, -1.1819432, 0.0448609, -2.9301040, -0.9612910, 0.6980560, -1.8484948, -0.8794564, -0.6786223, 0.1581767, 0.1375317, 0.1314209, 2.3444036, 1.6029342, -2.8400878, 1.1561869, 2.9171159, 2.4135232, 1.5075542, 1.1320685, -0.5064856, -1.4678970, 2.2886302, 1.3389820, 2.8791109, -2.9990327, -0.9727779, -1.1293601, -0.5565553, -1.8922157, -1.1486180, 0.1280838, -2.4063617, 0.4363001, 1.8407839, 0.0623114, 1.9006301, 2.6541438, -0.9666587, 1.9558349, -2.1466769, 2.5258323, -2.7064216, -1.0078697, 0.0972503, 2.1965265, -1.6650136, 1.0713067, 2.7244384, -0.0239241, -1.4176964, -1.5307467, -0.6815083, 1.9868009, 1.9384541, -2.2222969, -2.3594449, -0.7108697, -2.3041478, 2.8371039, 1.5034469, 2.4084996, 2.3496337, 0.5800164, 1.6029149, 0.6477948, 2.2794893, 1.4549921, 0.2358253, -2.6519530, 1.7865842, 0.7485075, 0.7219914, 0.8224096, 2.5169840, 0.4046851, 2.4150432, 2.7774971, -1.9893979, 2.5610111, 1.9568627, -2.1906926, 2.4437791, 0.3398526, -1.9971111, 1.3331908, 1.3366502, -1.6640590, 0.1541922, -1.3511698, -0.7559710, 2.3123246, 0.5964285, 2.8495858, -0.2675055, 0.9130170, -1.3038093, 1.8532567, 0.6015567, 1.5396335, -1.2245601, -2.2675414, -1.2598734, 0.8713270, -1.1092104, -0.8468686, 1.0034800, -1.5930650, -0.9039785, 1.7621119, -0.7921444, 0.5762513, 2.9613404, -2.2330469, 2.2239777, 0.2017585, 1.3712430, 0.0601386, 2.2101644, 2.7784161, 0.2273965, 1.0026569, -0.1511447, -2.7025221, -2.5021329, -2.9136918, -2.4059980, -0.8674049, -1.1181450, 1.5463757, 0.4721983, 1.8437893, 1.9628431, 1.8442487, 1.4583150, 1.9447717, 0.2692401, -1.1141738, 0.1936885, 2.8049695, -2.0893869, 1.0013960, -2.8819210, -0.8101856, -1.1556842, 0.2063261, -0.7058416, 1.4948662, -2.8777728, -0.2445889, -1.0679634, -2.8969254, -2.4999884, -1.0727212, 2.0008625, -2.6487970, -0.1455326, 2.2202447, 0.7238012, 0.1644317, 1.9650229, -1.5686900, 0.4907637, -2.4188214, -2.4423048, 2.6758256, -0.7006323, 2.0815592, 0.1908102, 1.9451768, 1.0664558, 2.9749635, 2.4418827, -2.3596827, -1.1685406, 0.7026694, -1.3133470, -1.6538908, -2.5877950, 1.3374262, -2.4947721, -2.2016080, 2.5367505, 1.3365001, 2.2332979, -0.4681284, 1.4224907, 2.0124960, 1.2643145, 2.8322120, -0.7603844, 1.9759344, 2.5049433, 0.3568433, 0.5046418, -2.0148691, 0.0783498, -0.9989950, 2.4288048, 2.6805458, 1.3921891, 1.8541908, -1.1322085, -2.8953986, -2.6653515, -2.2132848, 2.3927540, 1.8766861, 2.1394429, -2.3918123, -1.4434141, -2.5891833, -1.9859279, -0.4147315, 1.4258775, -1.7412499, -1.4038880, -0.7892727, 1.6019137, -2.5538856, -2.8000863, 1.2913798, -2.8160866, -2.2109570, -1.6859662, 2.9808178, 2.7991446, -0.8105781, 0.4024184, 0.5748475, 2.0064012, 1.8570438, -0.4964737, 0.9829818, 2.4031670, 0.2307517, -2.7855286, 0.1131501, 0.0689469, 2.6611622, -1.2936841, 2.7957905, 2.9595771, -2.6850132, -1.2931041, 2.0263037, 0.9315793, 2.1524555, 1.2427025, 0.9178514, -2.9044594, 1.1458232, -1.4179260, -2.1693960, -2.4075309, -0.2217481, -2.4123718, 0.9378804, -0.8461562, -0.1176234, 1.0551878, 1.6672317, 0.9086787, -2.1288690, 0.5356995, -0.1723102, -2.8177807, 1.9432006, -1.9231695, 1.1535202, -2.3289934, -1.1954392, 2.5514795, -1.5798375, 1.7355229, -0.9717965, -2.8332350, 1.5969503, 2.8662405, -1.3859814, -1.9042166, -2.7619679, -1.4217447, 0.8571960, -1.9262289, -0.4539641, -1.1867861, -0.7110415, 1.8485006, 0.0967604, -2.6863804, 0.1567643, 1.9300770, -2.8298082, -2.3665223, 1.2316671, -0.7798403, 2.3557780, -2.8283817, -1.8453802, 0.4999958, -0.1212104, -0.5836840, -1.4244176, 1.9684523, -0.6006388, -2.7847342, -1.9820542, -0.9300619, -0.3512381, -0.2427254, 1.8245204, 1.4717728, 1.0900468, 2.4330695, -0.4027966, 2.9076576, 0.1389746, -2.7568643, 1.9443199, -0.5612527, 1.9664390, 2.8892166, -2.5988985, 0.0276338, 1.9369831, -0.3916827, 1.0502736, 1.7531601, -1.9287048, 1.2150770, -1.3737767, -1.8664701, 1.8394620, 2.6446689, -0.6266738, 1.5494938, 0.0735751, 1.0331504, 0.9909551, -2.4778152, 0.9414086, -0.4146873, 1.4054984, 1.1804910, 2.0645974, -0.0945039, -0.5229170, 1.4095464, -0.4808584, 1.7576865, -2.8241118, -0.3964416, -0.0100525, -2.0714102, -0.4999668, -0.9648530, 0.9542874, -0.4956125, -1.8944908, 1.1449716, 2.4553697, 0.2899434, 0.7590899, 2.0549266, 0.8896686, 1.4611554, -1.5732205, 2.9368019, -1.6616264, 2.9702700, -0.5947345, -1.7335056, -1.2231479, -1.5250462, 2.0442651, -0.9485720, 0.4947795, -2.0630847, 1.6543401, -2.1504577, 1.9301274, 1.6289531, 2.3710380, 2.0931904, 1.9012275, 2.3154353, -1.7917307, 1.6497323, 2.5832783, 1.2192579, 1.4112977, 2.3318862, -2.7664505, 1.3596217, -2.1997426, -0.8944603, -1.9187457, 2.5807647, -0.3435832, 2.6564666, -0.9085469, -2.3637653, -2.4152136, 1.7411289, -0.2098545, -1.9381045, -1.7564107, 1.5859244, 1.2689313, -1.2725282, -1.9633896, -0.8221298, -1.3519394, -2.4670072, -0.1342302, 0.9067911, 0.7681947, 1.7568208, 0.7418147, -2.2915934, -1.3094740, -2.9041633, -0.8615687, 0.8316432, -2.8840405, 1.5208216, -0.0650652, -2.6278034, -0.1891730, -2.9975898, 0.4561515, -2.6782825, 1.2380775, 2.4959879, 1.4340504, -1.2531053, -0.2857239, -0.0297542, -1.8545757, -2.2358399, 1.9209761, 2.2578361, 2.9870241, 0.7113778, 1.7232219, 0.3435943, 0.9273232, -0.1629446, 2.6441357, 2.7309571, 0.3907827, -1.7036447, 2.2370898, 2.9023449, -2.0185947, -0.3379818, -2.6355685, -2.7084232, -1.0192767, 0.4783619, 0.2793264, -1.0605596, 1.7415567, -0.5320163, 1.2662667, -2.2058056, 1.6272680, -1.1352461, 2.3162938, 1.8337025, -2.5842385, 2.1055818, 0.9062107, -2.4067405, 1.3537672, -1.1653866, 2.1832775, 1.4171873, 2.5429260, -1.5022635, -0.6415177, -0.6940488, -0.5427436, 1.2202540, 1.0624286, -0.5663515, 1.9078589, -1.9688310, -2.8067301, 0.9455712, -1.5219181, -2.3934467, -1.6590911, 2.4750791, 1.0379790, -0.3523515, -0.9713846, -2.4951324, -1.3076749, 0.1624590, -1.6309914, -0.6556567, -2.1278697, 2.3827470, -0.6974015, 2.3263880, 0.6204501, -0.4442495, -2.9358908, 0.6158195, 2.8094546, 1.0322040, 1.2074609, 1.2319042, 1.7886505, 0.8644633, -0.1111528, -2.8547221, 2.8594324, -2.0691451, -0.1205691, 1.0929353, 0.5667916, -2.2711797, 2.6928191, 0.4816360, -0.9190635, -1.3500198, 2.3763000, 1.8443355, -0.3277826, -1.6989197, 2.1586755, -0.0816870, -1.3318819, 2.6130793, -2.2833754, -2.8996981, -2.9589714, -0.8713316, 2.7960791, -0.3252853, 0.7279752, -2.3111297, 1.8764362, -1.8069921, 0.1662807, 2.2140996, -1.2966107, 2.4675120, -0.3003752, 2.5054515, -0.1535400, -1.9301191, 0.3212296, -1.5259077, -2.6889680, -0.2955750, 0.1957438, 1.9816890, -1.7802980, 0.4444920, 2.9716527, 2.1098536, -1.2336314, 0.5313826, 2.9851955, -1.0439388, 1.2689216, 0.0923657, 0.6302680, 0.1521022, 1.8217356, -0.7744516, 0.1972817, -1.1803089, -0.6583296, 1.6797122, 2.1498977, -2.9455201, -2.7741093, 1.8546140, -1.1568670, -1.9506440, -1.1530780, 0.4886893, -0.6123114, -0.6670609, -2.1783698, 0.7011458, 1.7397908, -0.6028400, -2.8707296, 1.2155518, 0.3080017, -0.0114162, 2.2270849, 1.1076363, -1.3410047, 1.4625600, 0.3498712, -2.1632722, 2.0648997, -1.3626235, -0.8378344, 2.0816387, 1.6434224, -2.1987649, -2.7057182, 1.5196161, 2.2746137, -2.2332868, -2.2080967, 1.6593326, 1.9490996, 0.3490607, -1.9458467, 2.9447674, -0.6720046, -2.9147023, -2.2293491, 2.3246154, 2.2099504, -1.8731250, -1.2142976, 0.3050568, 1.2882323, -1.3380342, -1.5149851, 0.7835526, 2.4923613, -2.7750587, -2.5813610, 0.9325782, 0.2169591, -1.2668638, 0.5367069, -2.7711950, 2.4172189, -0.7046620, -2.4613199, 0.3217813, 2.4983133, 0.5728294, -0.2491716, -2.9135823, 1.4897410, 1.1677372, -1.8431406, 1.8749216, 1.8215466, 2.2320122, 1.5066070, 0.8120441, -2.0260641, 1.9611478, -2.5558942, -0.2675641, 2.0759875, -1.7840068, 1.2574455, 1.0346843, 2.6247657, -0.8165324, 0.7059279, 2.0144258, -0.3199139, -2.8949273, -0.2279426, -1.7406392, 0.5525624, -2.7317135, -2.5821404, -2.9027357, -0.1738188, -1.7971142, 0.4453376, -0.1635371, -2.2625403, -1.1884885, 0.5223974, 0.2093644, 0.2669993, 1.3667127, -0.4042958, -1.9141356, 0.2183450, 0.4099742, 0.9177399, 1.7252594, -1.5671473, -2.1057804, -1.1044032, -0.6383964, -1.7245748, 0.4405033, 2.2762208, 1.0734616, -0.5503442, -1.2440209, -2.9429006, 2.1150245, 0.4186177, -0.4522529, 2.0871342, 2.5826129, 1.3040903, 1.4532772, 1.2240798, 2.2726813, -1.8052528, -1.0809376, -2.0302163, 0.8697546, -1.5123862, -0.7009964, -0.4615629, -1.3026857, -1.5876839, 0.2475589, -1.8478794, 1.8911684, 2.2524428, -1.0652432, -1.7776209, 1.4241786, 1.1486429, -0.2296096, -2.0626586, 2.5104510, 0.9931582, 1.9858726, 2.3392785, 1.6319038, -2.7922218, 2.4118975, 2.8163235, 2.6115291, 2.9699124, 2.2142580, 1.6299426, -0.1192659, 0.4255255, -2.6753028, -1.4729919, 0.7961154, 1.6274480, 0.0740061, -0.8553317, -2.0620675, -1.9139055, -1.8596326, 2.4927596, -0.3923496, 0.8438519, -1.2692031, 0.4948120, 0.9839259, -1.3639838, -2.1822008, -0.9217124, 1.9445149, 2.0494097, -1.4829166, 0.4344227, 0.5197572, -0.6406347, 2.3655870, -1.2319096, -1.3070147, 2.5998868, -2.0267481, -2.0041843, -1.7961750, -0.9172319, 1.7086164, 0.1072215, 0.7321609, 2.3244316, -1.1405531, 1.2058596, 0.3654508, 2.3223165, 0.2337208, -1.1377241, -2.4082831, 2.5479789, 2.7700905, 1.4735067, 1.4487188, -0.6219324, -2.5100050, -2.9885489, -0.9361673, -2.5834981, -1.1703406, 1.7560932, 0.2145728, 0.0493131, -0.3947284, -0.7828327, -0.9829593, -1.5907749, 1.9443790, 0.5055910, -0.1364159, -1.4896622, 2.5475995, -2.9198976, -1.2760543, -0.6091050, -0.9088413, 2.5297358, 0.0865890, 2.6887338, -1.9699065, 1.8886529, 1.8704576, 1.0574723, 2.1784756, 2.0106160, 1.9395005, 0.1232729, 0.4564465, -2.5261567, 0.6432857, 2.8459252, -0.7376637, -0.3359882, -0.0565007, -0.9764024, 1.5025612, 0.3788087, -1.3870051, 0.6072691, 1.1190695, -2.8795421, -1.5366612, 0.7525938, 0.8214664, 1.6498288, 2.7634227, -1.4221412, -1.3394239, -2.3715841, 0.1236655, -2.5579599, -1.1385257, 0.0380517, 1.5278787, 0.5614509, -1.9870041, -1.6394684, -0.0547306, 1.4370022, -0.7179165, -2.8695628, 1.1896270, 1.1351775, 2.6197539, -0.0362031, -0.8215702, 0.9094319, 0.2991361, -1.5157274, 2.8037998, -2.6489147, -2.1076396, 2.6272552, -1.6625797, -1.9975139, -0.4670604, -0.4315071, 2.6186756, 0.7276883, 2.0571087, 2.8295514, 2.3289516, -1.8535367, 2.0529521, -1.2113356, -0.3684771, -1.4563413, -1.6963880, -2.2735810, 2.8061204, -2.6669562, 0.9795710, 2.0414215, -2.0335257, 1.7249085, -1.6256522, -2.7671742, -1.3185195, -2.0770245, -2.5941552, 0.0872069, 1.0467152, -1.0564255, -1.9685888, 2.2961557, -0.4400046, 0.1029708, -2.4608604, -2.1662958, 2.4128527, -1.8932100, -2.4332663, 2.1746559, -1.8760249, 2.1204558, -2.5557433, -2.2948185, 1.8423283, -0.5267944, -1.0865120, -0.6380755, -2.4056083, -2.3531727, 2.2389998, -2.8615296, 2.0556632, -1.3198462, -2.3350872, -0.3384871, 0.6137025, -2.9829225, 1.2123900, 0.2748409, 2.4206402, -2.0140916, 2.3010346, 2.7595265, -1.8034073, -1.9370535, -0.2368420, -0.4932976, -1.5002207, 2.3553688, -1.4537485, -2.9394147, 0.1413182, -0.9860493, 2.9415674, 2.7014428, -2.7390459, -1.5860119, 1.7954677, -2.0601402, 1.0214331, -2.2942722, 1.4179780, 1.2363904, -0.4722549, 1.4876522, 2.9984467, -0.8376742, -2.4135981, 1.0441584, 2.8107191, -2.6057353, -1.5758426, 1.2217885, 0.5284420, 1.1037361, -1.9534363, -1.9705591, -2.5718748, -1.3669759, 2.1369575, -2.1018852, 2.9973947, 2.0408508, 1.4770036, -0.7987212, -0.1301664, -2.7481288, -2.7384263, 1.2843399, -0.6770837, 2.1269483, 1.1205382, -1.7941849, -2.9232718, -2.9547399, -1.7345619, 1.8812156, -0.1932412, 2.4746867, 2.3360891, -1.3524425, -0.2055749, 0.4744215, -0.8746264, 0.1657838, -0.1675483, -2.1513608, 0.1366231, 1.0997731, -0.8799453, 0.7977385, 2.5769027, 0.6384327, -2.8511719, 2.6733198, -1.4272978, 2.6250150, 1.1173937, 1.9242434, 2.8883310, 2.7518507, -0.5327570, -1.0179736, 1.7374323, 1.2920684, -2.5856075, 1.9607971, -2.6961675, -2.2340458, -1.7885914, -2.9371562, -2.9824638, 0.7211701, -2.5556244, 1.7885009, 1.8406392, 2.8490077, -1.8778296, -2.1632928, -2.3411964, -0.3549621, -0.9664225, 2.1537495, -2.8646982, 0.5576591, -1.0833487, -1.0120086, 2.3985866, 2.5675574, -2.6127118, -2.8119984, 1.7168299, -2.4151002, 2.6976172, -2.9033222, 0.6210693, -2.5173000, 1.1696758, 2.6341833, 1.7964597, 0.1189138, -1.6117093, -1.8061677, -2.8835053, -2.6212343, 1.3216061, 0.3053065, -2.7802989, 2.3072443, -1.5819037, 1.4729558, -0.9055460, 2.7831603, 0.2805882, 0.5312444, 1.5031648, -1.1994395, 2.1699708, -0.6502802, 2.5476584, -0.1203106, 2.0370550, -1.8118306, 2.2926617, -0.1674348, -2.5844001, 2.8794346, 1.0947871, -1.4925987, 0.7968500, 0.4269043, -0.0021779, 2.9628030, 2.7683208, 1.0658141, 0.2068065, 0.8475730, 2.0120073, 2.5881325, -0.0974500, -2.4556339, -1.5954025, -0.4639675, 1.9369112, 1.7674934, -0.6670460, -0.7490566, -2.3154713, -0.2979497, 0.2633435, 1.9589228, -0.4814294, 2.7527862, 1.7785361, -0.9635706, -0.2142536, 0.6939435, 1.8346836, 0.7357150, 0.3137520, 2.0397089, -2.2017772, -0.6293449, 2.8396616, -0.2411100, 1.8818074, -0.3114219, -2.9093264, -2.1145643, 0.8276870, -2.0590954, 2.2222879, -2.7449154, 2.3391556, 1.8064191, 0.2878009, 0.0505901, -0.6176663, -0.3635876, -2.6063475, 0.3111487, 2.0894362, -2.3779299, 1.6395500, -0.7055607, -0.4347288, 2.7382813, 0.4400229, -2.0431870, -2.5986720, 0.7653862, 0.1704355, 1.4921829, -0.9709304, -2.0896703, 1.9222186, -1.6816066, -0.0554982, 1.4926263, 1.1964506, -1.9544337, -1.4860663, 2.1342098, 1.5675222, -2.6762343, -2.5071386, 2.9919429, -2.8241980, 2.4852741, -0.7818139, 0.7623761, -2.4900820, 0.7055096, 2.7214221, 1.0319331, 0.7696510, -2.7738648, -2.1153144, 2.6830560, 0.3908663, 0.8111929, 0.8002455, 0.2505208, -0.3176185, 0.5661428, -1.6464027, 0.2261498, -0.6521966, 0.0033654, -1.4520710, 2.3951754, 1.4233837, -1.7413166, -2.1852894, -1.2826303, 0.9150687, 0.5253614, -1.9686453, 2.2720309, -1.4798541, 0.5099374, -0.1167664, -1.5252278, 2.7682805, -1.9340241, 2.7396781, -2.2724923, 2.1335230, -1.1198255, 2.5096704, 2.6717960, 0.8339812, 0.4756174, -0.6992569, 2.0414848, -1.0503495, 2.6843217, 1.7253941, -2.5993834, 0.7806892, -1.5986134, 1.2905872, -2.1634159, 2.6071157, 1.9212036, -1.5892957, -2.0262513, 0.7265411, 0.1145224, -1.3373205, 0.6821852, 1.7670741, -1.4222790, 2.2067335, 1.5131488, 1.6626174, 1.4326072, -1.1987955, -2.3912152, -0.1736365, 0.4905701, -1.2838712, 2.4556928, -1.0957366, 0.3303268, -0.9658985, -1.8478107, 2.6042505, 1.6228499, 1.7742812, 1.6238811, 0.2763472, 2.9583530, 2.5610072, -1.8642833, 1.5805283, 2.7585425, -0.4782475, 0.1132706, 1.7917236, -1.7963705, -2.3302647, -2.4841882, 1.0922242, 2.6939962, -0.1722397, -2.0268667, 2.2425456, -2.9343930, -1.7465186, 1.1376526, 2.4884983, -1.9998624, -1.1599949, 1.9942312, 2.4682658, -1.3553675, 1.1896391, 2.5058415, 0.4419614, -1.9258681, -0.8388414, -2.3124579, -0.3666370, 0.8644476, -2.5536347, -0.3451603, -1.7805529, 1.9814342, 0.4222204, -0.9595745, 1.8066377, 0.8501171, -2.6579053, 0.3797355, 2.0244854, 0.7383596, -0.1410795, -0.7204138, -2.8847948, 0.2162639, -2.3660260, -0.5745967, 0.0647568, 0.5258108, -0.6554541, 1.7625407, 0.0877316, 0.6454362, 2.2215048, -2.1179414, 2.1549047, 2.3521624, 0.2771448, -2.7489398, -2.9515141, 1.8838575, -2.3238797, -1.4989653, -1.0816376, -2.5061178, -2.5149767, -2.2494947, 1.2590269, 2.4980556, 1.4045319, -0.5090745, -2.1497761, 1.7552358, -2.2273017, -1.7790727, 2.5950440, -0.7588872, -1.6150220, -0.7793858, -1.9255352, 0.9157256, 0.7778540, -0.7330852, 2.3978169, 1.2191753, -0.0699772, -0.5106853, -1.6627672, 0.2854112, 1.8387018, 1.6959513, 1.4414453, 2.5824540, -0.1309801, 1.1646637, -2.8680072, -0.1028627, -1.0474153, 1.0589897, 1.6425075, 0.7393063, 2.1582168, -1.2387909, 2.3122597, -2.0170995, -1.6660732, 1.1285682, 2.8302578, -1.2893007, -2.6458561, -1.9487873, -0.9764827, 1.3997158, -0.6430854, 0.1954877, -0.6922585, 0.0537666, 1.6483464, 1.5670097, 0.9843719, 2.9123453, -0.5010517, -1.5782922, -1.9182365, -0.7396289, -0.6009301, 2.4050151, -0.7230319, 1.9113267, -2.9846422, 1.9829146, -0.8320269, -0.5115907, -0.3920738, -2.5383914, 2.0159650, -1.6431232, 1.1776784, 0.9030317, 0.0045884, 2.2153099, -0.1320079, 2.5744253, -1.0226142, -1.6449557, -1.2032224, 2.2722968, 0.0627049, -0.4289228, 1.0946761, -2.9065164, 2.7910944, -1.3791682, 2.4262208, 2.5055603, -2.1177706, 2.1605181, 1.3960859, 2.6120725, 1.5405531, -0.9094227, 1.1717347, 0.5650308, 0.2330681, 0.8399154, -0.0335606, 0.0283195, 1.7264228, -1.7382459, 2.5355245, 0.5053993, -0.3936678, -0.2592107, -0.9273910, -1.8856868, -0.5731207, 0.2239504, 2.6999986, -2.9766651, -2.3304416, -1.4987850, -0.7608706, 0.1710580, -1.2839339, 0.7991638, -1.1325126, -0.1303038, -1.8587785, 1.6897318, -0.8002624, -0.4782266, 0.9863480, -0.9930927, -2.1511240, 2.2001628, -2.2911738, -1.5422669, 0.2960820, 2.9318757, -2.4056098, 1.6454914, 1.4238039, 2.8656887, 0.2858998, -0.3873639, -1.6227329, 0.4839268, -0.1960562, 2.6989245, -1.2597767, -1.2222372, -2.9176837, -2.4136528, -2.1218078, -1.4342398, 1.8076489, 1.1325593, 2.1665430, 1.0374454, -0.8277341, 0.9004040, -2.8552974, 2.2246879, 1.0038141, 1.3710962, -1.2063226, 0.7115140, 1.6492871, -2.8365560, 0.3741179, -1.2184286, 2.9752362, -1.1534710, 2.4660195, -0.5926808, -0.3045739, 2.2569941, -2.9226311, 2.7002166, -1.2087629, 2.7654322, -2.9428146, -1.7773958, -0.6687404, -0.7511282, -0.0512626, -2.9803172, 2.5440447, 2.1545139, 1.9877289, 2.6189632, -1.8336718, 1.6383965, 0.6509851, 2.3947896, -2.7767276, -2.2975965, -0.5571612, -0.2503024, 2.9520396, -1.1230466, 0.1008542, 1.9125704, -2.5164831, 0.0230511, -2.5787483, -2.2697826, 1.2145138, -1.8529628, 0.6324264, 2.8998598, -0.3379567, -2.2605740, 0.5203199, -0.7662181, -1.9289942, -2.4102796, 1.4628472, 0.6499326, -2.1896977, 2.5117385, 1.9538500, 0.7061858, -2.9990367, -1.2864451, 0.9234093, 0.8479439, -1.5153478, -2.0461048, -2.8234358, 1.6782149, 0.1121689, -1.8350652, 0.9130173, -2.1153918, -2.7160704, -2.8871187, -1.7879538, 1.0681458, -1.6430170, 0.0378467, 0.9261964, 1.7191195, 0.8087080, -2.3199122, -0.7230456, -1.5640887, 0.4028205, 2.2439474, -2.5808606, 0.4997607, -0.8368311, 1.8425746, -0.5435689, -1.0715483, -2.4694077, -2.0392261, -1.8364282, -1.2467503, 2.0772525, 2.0885065, -2.9842533, 0.0735410, -1.8486499, 0.7407991, 1.5862519, 0.6257154, 2.3662930, 0.2385068, -1.6026994, 0.8043314, 2.8990508, -2.6124941, -1.2252659, -0.8453659, -1.2712221, -1.4332534, -0.3839940, -0.2833051, 2.9392893, 1.8242194, 0.3488436, -0.5158334, 1.7239477, -0.4713857, 1.5907595, 0.4606923, -1.5792053, 0.5149298, 0.4909076, -1.5629317, 1.7935706, 0.1298317, 1.2965691, 2.2286807, 1.0843116, -2.2554043, -1.6335147, -1.7600546, -2.3498448, -0.3197840, -1.0202439, -1.8977156, 1.6947917, 2.7335045, -2.0617959, -2.3877442, -0.5658121, -0.8489251, -2.8269870, -2.3689773, 0.5934419, -1.8273538, -1.9043678, 1.7689259, 1.4356529, 2.3237876, -2.7222270, -1.7987001, -0.6615503, 0.5797769, 0.5104594, 2.3565847, -0.1732453, 1.6489884, 1.9455803, 0.1705114, 2.4472897, -2.3356494, -1.0543600, 0.8826526, -1.3021243, -2.3760779, -1.9263480, -2.8719494, -2.8269500, -2.7369948, 1.7965395, -2.2117849, -2.6053038, -2.2044229, -1.1421135, 0.4467279, -0.6462072, -1.3795599, -1.4928610, -2.9442969, -1.9804527, 2.3348863, -0.3935945, -2.3769456, 1.4046082, -0.2620207, 1.1849497, -0.4190337, 2.6653776, 1.9582333, -0.6551991, -1.1061484, 0.9322603, -0.9391485, -2.7753320, 2.5713989, -2.7252632, -0.8773454, -1.9385097, 2.2465426, -1.1058288, 2.4638689, -2.4264060, 1.8328402, 1.0340660, -1.5501588, -0.8855823, -0.0686690, -2.3748005, -1.0733233, 1.5341866, -0.6816694, 0.7254371, -0.2553383, -2.5248459, -2.8307591, 2.0812425, 2.0653225, -0.7631544, 2.7220023, 2.5167757, -1.5189002, -1.2490956, 0.2503877, -1.3911689, -0.0611133, 0.8749186, -0.0361843, -2.5876892, 0.5525846, -1.6218174, -2.2479038, -0.5315124, 1.3081987, -0.6091996, -2.4715295, 1.2351183, 2.0879709, 2.5692245, -0.4019676, 2.9533557, 2.9342209, -1.1682357, -2.5785822, 2.9549707, 0.0490608, -0.0160013, -2.4307684, 0.2890703, -2.2460507, 1.5100827, 0.6329676, -0.9698253, 1.2186022, -2.1639148, -1.5212618, 0.7230886, 1.0044733, -1.0611762, -2.8240093, -0.4443458, -0.5742865, 2.0609146, 1.0785600, -1.1315282, 2.2875879, -1.7195962, 1.6522241, 2.7026249, 0.9551203, 0.4468619, 0.4060567, -2.6887149, 2.9759668, -2.0125402, -0.1209857, 0.7586776, 2.3677110, 1.0759299, 2.4904592, -1.9442604, 0.2491843, -2.6134877, -0.5970973, -0.0492762, -0.4628646, -0.1720775, 0.1091746, -1.6567423, 0.3969552, -0.3900869, 1.3849734, 0.0061245, -1.9941746, -1.8905827, -0.2920612, -1.1758580, -1.4790636, 0.2200756, -0.1499835, 0.0710421, 1.7811435, 0.6053707, 0.3455518, 1.6601846, -0.3478340, 1.2109605, -0.9152858, 0.8394999, -0.5699171, -2.4420733, 1.3955426, -2.6635962, -0.8885802, -0.4328569, 1.9790669, 2.6845549, -2.2328747, -0.3989024, 0.0809444, -1.6973512, -1.8550108, -0.9776302, -2.3468466, -0.2748405, 2.2068024, -1.3648404, -2.5564387, -0.6450383, -0.8147452, 2.6985462, 1.3253641, 0.9286326, -0.8660231, -0.1863761, -0.1619888, -2.2873280, 1.5484511, 2.8052243, 2.6233191, -2.6347413, 2.5943041, -2.1253839, -1.5330329, -2.7699105, -2.7721166, -2.2000522, 1.6178803, 2.2249443, 1.2373182, 1.8636238, -1.3913594, 2.5014740, -1.6500907, 0.1125542, 2.7295381, -2.0509357, 1.9539632, -1.8249491, -0.2727357, 1.2901407, -0.1706969, 0.6288947, 2.9841251, -0.8412379, -1.8740278, -0.8962678, -1.3000556, 0.8666047, 1.2667804, 2.5785196, 0.0033394, -1.0685235, 1.4845530, 1.3048864, 1.5464746, 2.4378493, 0.3599194, -0.5992526, -1.5133375, -0.1321313, -0.4315924, 1.5955667, -1.3710371, -1.9236157, 0.2008691, -0.5264382, 2.0305645, -2.2882134, 1.1879073, 0.7059526, 0.9690112, 1.6219567, 2.9551418, -1.3387821, 1.7333809, -0.6037193, -0.0624041, 0.7890569, -0.1601556, 0.9172313, 2.4472634, 1.1586377, 2.3722551, -1.7589119, 1.8200348, -0.6250559, -2.1306361, 2.6075889, -0.6576097, -0.9383336, 0.6671527, -1.9459892, 1.8185712, -2.2948370, 1.8593325, 0.2074865, 2.8331754, 0.3019502, 0.5420654, -0.0378859, -1.8091190, 2.7689125, 0.2558574, 1.2088823, -0.1610995, 1.4123210, -2.8010245, -1.3285136, 2.2970950, -2.4062790, 1.4230136, -0.0372803, 1.3591109, 0.7431981, -0.2291804, 0.7996581, 1.1367367, -1.3334636, 2.1584375, 0.9675677, -1.8211412, -2.0251265, -2.9327024, -1.7775001, 2.4448113, 0.4844407, -2.8951697, -0.3513374, 0.2545000, -2.4865677, -2.2832573, 1.5595762, 2.9955513, -0.9458991, 1.6430514, -2.5881512, 0.5986014, 0.8666653, -2.7780706, 1.4398401, 2.9549748, -2.9650817, -2.0075120, -1.5438715, 1.8671510, -1.3830760, 1.5271402, 2.3506791, 1.6858140, -0.6530256, -2.7588546, -0.1376826, -2.9864634, 2.4907296, -2.4044673, -2.7827465, 2.6855313, -1.1338435, -0.2710101, -1.9754660, -1.4711006, 1.0764572, 2.4492420, -1.6989698, -0.3837878, 0.9326389, 2.5571309, -1.0357715, -0.7615785, -1.0398625, -1.2055175, 1.1292209, -0.6090180, -1.8900193, -1.2604224, -0.6654873, -2.0814913, -2.4535350, 2.8764464, -2.5055788, -1.4851071, -1.2124818, 1.2843701, -1.1252210, -2.5844892, 0.3268405, -0.3577003, -2.2368378, -1.0018747, -1.6348277, 0.7458628, -1.3034273, 2.4561876, 0.0072334, -1.8272728, 2.2754477, 2.5557031, -1.8866244, -0.6545107, 2.8739453, -0.8368037, 2.4020478, 1.3719145, 2.1789721, 1.4135459, 1.8816382, -2.6460301, -2.5202059, -1.4222883, -2.7520458, 2.5552235, -1.9394228, 0.1074765, 1.8612872, 0.8670754, -1.5043098, 0.8813025, 2.5358419, 1.9867205, 1.2085742, 1.7528566, 0.0596301, -0.5995150, 0.4727775, -2.8602574, 0.7101019, 1.7273714, 0.8666942, 0.6807091, -0.3583623, 2.0687235, 2.7711887, 1.1327389, -0.3778020, -2.2451612, 2.2350846, 1.5491663, 1.4532563, 1.2127786, 0.8418527, 2.6101150, 2.7367225, -2.3923187, 0.3985145, -1.8238132, -1.5379171, -2.3902486, -1.2914220, -2.6977872, -0.7384476, -1.0496028, 1.2923524, 1.3956059, -1.4761863, 1.2097430, -1.1190730, -0.5415709, 1.6595996, -0.5543355, -2.3464852, -1.3794360, -0.9360298, -2.2385964, 1.0088166, 1.9726423, 0.9725690, -1.9998057, -1.1749931, 1.4858852, -0.1039561, 2.0758910, 1.2204588, 2.4963570, 0.8295068, -0.4745570, 1.2016148, -1.1956714, -2.8196039, -2.4951124, 2.8302958, 2.6192827, -1.3653963, 0.0183039, 2.4081423, -2.2462548, -2.0636296, 2.4540888, -0.5486021, 2.3941076, -0.4291531, -1.5876420, -2.6297766, 2.5911487, -0.4423385, -0.1181789, -1.4949818, -2.6187786, 2.5240007, 0.8802138, 1.5463030, 0.5642550, 2.3349616, -0.6249198, -2.0257687, -2.6515975, -2.9214429, -0.7778932, 1.9091932, -1.5667201, -1.7241212, -2.3304837, 1.2728336, 1.8983501, 1.9837205, -0.8894651, 0.2126234, -0.7130042, 2.5374117, -2.3190181, 2.1912764, 0.0434800, 0.4877658, 0.5028887, -2.9420027, 0.8224278, 2.8839432, 0.4608162, -0.3191136, -0.7320917, 2.1638883, -1.3303076, -0.1838740, 0.7342084, -2.4698137, -2.2569477, 0.2741757, -1.4233093, -1.7249013, -2.6077124, -0.1445159, -2.6521869, 2.2334723, -0.1290918, -2.1476020, -0.4706794, -1.3926768, -0.6351531, -2.1431413, -0.3928996, 0.6923323, -0.2006472, -0.9676461, -0.7035549, -0.5926451, -1.7494722, -0.4851778, 1.1186055, -1.0453773, -2.7543492, 2.5345241, -1.7150526, -2.3299854, -1.0454469, 0.7505579, 1.2705588, -0.9896628, 0.7009928, -2.4286781, 0.3868538, -0.5813335, 2.9367950, 2.8624624, -1.8531660, 2.4643859, -1.6345406, -2.8873474, -1.5750397, 1.8024490, -2.7020222, -0.0573321, -0.3416733, 1.8449356, -1.3923732, 1.3427675, 0.0999631, 0.8566921, -2.1702058, -1.1909378, 0.3761895, 1.2618387, -1.8651424, 2.1235096, -1.3898390, -2.1174312, -0.8506336, -0.1363864, -2.9496585, -0.8393277, 1.1419720, -2.9557563, -2.2502587, -1.6352461, 2.3246802, -0.5754469, 0.7917193, -0.9616588, -0.7078651, -0.5080451, -1.2471047, 2.4831963, -2.2465443, -2.1624357, 1.6162737, -1.1490719, 0.7667104, -0.0737654, 0.9492157, -2.3863431, -0.0117172, 2.4291044, 0.1652851, 1.0249889, 1.4996112, 0.7334290, 2.4971879, 0.7226641, 1.1489290, 0.1105860, -1.8446715, -0.0430896, -0.8604606, 2.5994797, 2.6949439, -1.7140735, 2.0114400, 0.3066455, 0.2712647, 2.0971424, -2.7859992, -0.4191172, 0.9092659, 2.1039389, -2.0720134, 1.9327156, -2.8352763, -0.2243825, -1.6883387, 1.7780247, -2.2422968, -0.9295672, 0.3971709, -1.1127891, 1.1828294, -2.9388748, 1.5626510, -1.6014486, -1.9765473, -1.6353552, -2.9844019, -2.7648776, 1.8803940, 0.0934908, 1.6393573, -2.0562353, -1.7563264, -1.8073598, 1.0480139, 1.0299923, 1.0315811, -1.3255473, -1.9488219, 0.4581183, -0.7119820, -0.9454119, -0.2053760, -0.7981751, 1.2156009, -2.8312420, -0.1191850, -1.5934823, 0.4339245, -0.5667886, -2.7531066, 0.6168024, 2.0356641, -1.0914795, 0.3364086, 2.3990753, 0.2825325, 0.9491197, -1.5449947, -0.5514503, 0.2112812, -1.5409094, -0.5777355, 2.2525793, -0.4141943, 1.8770764, 0.6103372, 0.4773493, 1.8311157, 1.3982844, -1.7452546, 2.1097550, -0.7444452, 0.6265396, 2.7278234, 2.4830765, 0.8170471, -1.3686222, 0.7300142, -0.8683378, -0.3895906, -2.1397437, 0.4612525, -2.7116841, 1.1126187, -2.7473962, -1.1772868, 0.3731675, -1.2450285, -2.1740504, -1.4195262, 0.1314615, -0.2509814, -1.6566169, 0.8932708, -1.0404423, -2.6973108, 1.7978155, -2.3119986, 2.6669974, 0.6520150, 1.7452582, -1.4350827, -2.2630788, -0.1839496, 1.6640936, -2.0894682, -1.6755804, -1.5515571, -1.2920254, 2.4908404, 0.5882049, -1.0525048, -0.1877540, -1.6910346, -1.3975167, -0.9648959, -1.4739095, -1.0079309, 2.9968437, -1.8200954, -1.7476173, -2.9646096, 1.0612751, 2.7477197, -1.4820926, -0.5784666, -0.7753818, -0.7995496, 1.1239214, -0.6480343, 0.8692727, -0.7321448, -0.9771900, -2.0374463, -2.1481084, -2.4843250, -0.5828665, 2.2852848, 1.6319564, -1.6371496, -2.0704524, -0.8563426, -2.4551324, 1.2871068, 0.7539484, 1.5004335, 0.6548880, -2.8140213, 1.6766018, -1.9025084, 0.5992198, 2.8668265, 1.6881722, -2.4663785, 0.6002124, -1.3838194, 1.0746494, -0.0400969, -0.2621395, 1.6864354, 2.6847226, 2.0006202, 2.7705150, 1.2687912, 0.9987735, 0.3516681, -1.7929669, 0.2932294, -1.4618415, 1.3229995, 0.9755869, 2.2967250, -0.4642916, -2.7999389, -0.0286353, -0.5808914, -0.2816400, -1.7544928, -2.2637507, 2.2894217, -2.7524994, -0.3265397, -0.4781458, -1.0214002, 2.4955358, 0.5872841, -1.3462596, 2.6327391, 0.9665605, -0.1787750, 1.9357173, 1.8538125, -1.7678082, 0.1042085, -0.8002423, -1.5217816, -0.2951520, -0.7795898, -0.8647668, 0.8333569, -2.8281256, 0.8056571, 1.4662890, 2.9619316, -0.2877662, -0.0050215, 1.0173443, -1.2239311, -1.1986691, 0.3623767, 1.8235330, -0.3540745, 2.7228601, -2.0454350, 2.5487395, 0.7126852, 0.7371348, -0.1691690, -2.2806778, 2.5771682, -2.2917664, -0.3301861, 1.6745946, 2.7711583, 1.9073308, -0.2596763, -2.7264305, 2.1614367, 1.6125989, 0.6126085, 1.3805340, 2.1912454, 2.3125690, -0.4194701, -2.8037022, 2.5901651, 0.7365711, -0.0949472, -0.5029826, 0.8775379, 1.1302814, 0.9829539, -1.7919900, 1.4777726, -1.1568396, 1.1889161, -0.7791800, 0.8497589, 1.5260805, -1.2722087, -0.1592336, 0.2665840, 2.9852199, 1.1495114, -2.0388222, 1.6388730, -0.0194914, 1.7525842, -2.6188986, 0.9538731, -1.8721631, -0.3747809, 2.3972933, -2.9628046, -0.0355258, 2.5352492, -1.7401162, -2.5413747, 1.6706722, 0.6803812, -0.5099698, 0.1179392, -1.1036000, -1.7217572, 1.0834010, -0.0158324, -2.9351787, 0.4970714, -2.3950087, -1.3407340, -2.4520535, -0.4775551, 0.3461324, -1.3358843, 1.6708218, 1.9871307, -2.0580719, -2.6589210, 1.6689634, 0.7688964, 2.6687795, 2.6902333, -2.0237888, 0.0717514, -0.1093135, 2.7336464, -2.9783101, -0.2641672, 0.6285615, 2.0429029, -2.7440505, -2.3813092, 0.3486140, 2.6679089, -0.8118718, -0.1815327, -2.7750626, 1.7852992, -2.6064140, 0.0185231, 0.0701162, 2.7634636, 2.1006630, 0.9745345, -1.8563658, -0.8248182, -2.7631863, -0.2107763, 2.1435353, -0.8234676, 0.6077797, -0.7557247, 0.9771295, -2.6281038, -1.8339702, -1.8821581, 0.1007531, 0.3829493, 2.5632435, -1.8799393, -1.8985408, 1.3994997, -1.1544050, -1.6952809, 1.8833231, 2.1815703, 1.8797908, -2.4366903, 1.8891488, 2.2719499, -0.3911267, -0.9888723, -2.8537969, 0.2836601, 1.2942488, 2.4755846, -0.9454658, 2.7541055, -2.0956984, -2.2370312, 1.1851108, 1.3599030, -1.3904059, -0.3961502, -1.5357691, -0.9109749, 2.8203860, -1.6809221, -1.9779585, 0.3017119, -0.0420821, -0.0294134, 1.6814209, 0.1162721, 0.2768561, 1.2328730, 0.0677898, -2.4803390, 0.3641549, -0.6803539, 2.3854146, -0.7769522, 1.8980052, -2.1756524, 1.8600867, 1.4056884, 2.3612452, 2.5029753, 2.0508822, 0.3131830, 0.7196771, -1.0481548, -1.6470017, -0.0509759, -2.7100037, -1.8003054, -1.7570416, 1.9413557, 0.8769556, 1.8482556, 1.5657968, -1.1105239, -0.9183746, -0.2924849, 0.9004381, 0.3418586, -0.5824477, -1.9498647, 2.9972490, 2.6670470, -0.6445060, -1.3707071, -1.9803849, -2.7325809, -0.5925820, -1.7424852, -0.3530136, 0.0159959, 0.0959464, 1.1765450, 0.9115742, 1.8790947, 1.2903454, 0.6553803, 1.3055043, 0.1956665, 1.0623634, -1.0449645, -1.0075189, -0.9984121, -2.6162115, -0.1277337, 1.1683758, -0.5953044, -2.8955899, 2.7194936, -0.2135879, -2.2321173, -1.7133267, -1.1251873, -0.8823082, -2.6041706, 0.3668257, 1.7445272, 0.8060610, 2.3072275, -1.3103072, -1.4333589, 2.5212072, -1.9742188, -2.8994047, -2.4255500, 1.1724096, 2.7634701, -1.3108700, -2.4148362, 0.5692289, -1.4233680, 2.4216471, 2.0237752, -2.5735734, -2.4598069, 1.8577601, -2.2709206, 1.7681218, -2.3072328, 0.9238703, 0.6574987, -1.7237567, -0.5031997, 0.5462858, 0.6021714, 0.8350926, -0.9357011, -0.4472976, 0.0120191, -1.5517098, 0.7516248, 1.3259842, -1.6552373, 2.9850645, -1.2677839, 2.7594507, 2.4923996, -0.0609771, -0.9891339, 2.4244492, -2.5288860, -2.6512858, 2.2062122, 2.9304262, -1.6424445, -0.7302796, 1.7216658, -2.9876548, -1.1723967, -1.9025690, -2.4900921, 0.1698577, 1.2581077, 1.0020883, 2.3104727, 1.6984156, 2.0176086, -0.2463337, -0.3685204, 0.5782550, -0.5757428, 2.7563023, 2.2726782, 0.5164129, -2.4961256, 1.3677865, 1.1692034, 0.3976342, -1.6149413, -0.2671664, -0.6478929, -2.5634043, 2.8598211, 2.9618252, -1.4821138, -2.0278359, -1.2610234, -1.3645501, 0.9720717, 0.8891347, 1.1636114, -1.1914794, -2.2301010, -1.2660120, 2.3670377, -0.9513956, 2.6188917, 1.0117444, 1.6092416, 0.7488641, 1.9249933, 0.0138285, 0.8900448, -0.1972414, -0.3514796, -1.6355637, 0.0812123, -2.2224018, 0.6175627, 0.0144496, 1.0863286, -0.8013766, -1.5613009, 0.8612201, -2.5279553, 1.3491592, 2.7859394, -0.3289700, 0.3829614, -0.1112770, -1.0431645, 1.8858598, 2.0750578, 1.9879012, 0.9211817, -1.3467241, 2.0503840, 1.1498697, 2.5917361, -0.5533701, -1.3413369, 0.2068209, -1.9828231, 0.8454753, 1.3708946, 1.9656843, -0.1177131, -1.6507641, 2.2724624, 2.1240240, -2.4415151, 2.8674729, -2.7226795, -1.5665694, 0.6744265, 0.4730840, -2.9545417, -1.0385807, -1.4467403, -0.4796573, -0.7091410, 0.4710779, -2.1475541, -2.8285875, 2.0874411, -0.7986251, 1.3804462, -1.5807558, -0.1480223, -1.5857401, 0.6082892, 2.6296299, 2.2550210, -2.0418336, -1.4768779, 1.4488425, 2.1391564, 1.5808504, -0.5184449, 1.3759940, -1.6313000, 1.9875814, -0.4022471, -2.4558636, 1.8025681, 0.4600112, 1.0081443, 0.6845191, 2.8119298, 1.4984881, -0.3810164, -1.5401851, -1.7139775, -1.0535924, -1.3770742, 1.4327816, 2.3177771, 0.2631205, 1.7509393, -0.8054755, 0.1846938, 0.8068449, -1.6939586, 0.0598269, 1.4222420, -1.3811323, 0.2609737, -0.3343638, 0.1596810, -1.8329229, -2.4540247, 0.1270381, 1.3965956, -2.4900475, -0.1406202, -0.8600071, 2.3013231, -1.0041229, 1.4319667, -2.8963529, 1.6531618, 1.0882376, 0.5946728, -0.6173265, 1.9245790, -1.5026098, 0.8033517, 2.7749949, -0.8258282, -2.0745595, -1.2348291, 2.8594638, -0.8049649, 2.0587227, -2.1602186, 1.6009460, -0.0227737, 1.2642943, -1.3400962, 2.4587423, 1.6937931, 0.0845069, -2.3405167, -2.5920035, -0.2982000, -1.9516784, -0.4250094, 0.7684446, -2.6427144, 2.1175473, -2.8353371, 0.7373804, 2.4185654, 1.2581669, -2.5436474, 0.2485767, -1.8701859, -2.6694787, -0.6400924, 2.6082479, -0.4873149, -2.2741677, -1.9729957, 1.3155876, -2.9798507, 0.9073137, -1.1712915, -2.7371301, 2.0313561, -0.8558014, -0.4016268, 1.2598113, -2.9238062, -0.3366974, 2.8415050, 2.2780693, -0.3892388, 0.4811362, -1.6535577, -0.4108041, -2.3813679, -0.1585306, 0.6483239, -1.4225788, 1.9625759, 0.3199607, -2.3675731, 2.6565770, -0.4265498, 0.5881232, 1.4629912, -1.3248964, -1.8527488, -0.1732675, -0.2000489, -2.4266307, -1.1486308, -2.6421217, -0.1352325, 1.2830944, 0.3436763, -1.1943372, -0.6178320, -1.7585969, 0.3310265, -1.0278677, -0.6459233, -0.6678994, -0.3882910, 1.2132411, 1.9787623, 0.4701074, -2.3433816, 0.7301065, -0.1808000, -1.3519672, 2.2477145, 0.1077421, -2.5811603, -1.0035610, 0.3600608, -2.8791340, 2.0014165, -1.8927848, 2.0329194, -0.2236753, 1.8061481, 1.6733149, -1.2286200, -2.1319335, -2.8261295, 1.5305991, -0.1322415, -0.3308702, 2.1005765, -2.1301660, -2.3365810, 1.6133430, -1.7269183, 1.1839859, -0.2915528, -0.8448710, 1.4563147, 0.9635714, -1.6498778, -2.5909279, 0.3479957, -1.5447094, -2.9121542, 1.1552517, -0.4350155, -0.2512793, 0.5826840, -0.2909766, 1.6861775, -0.5764945, 1.9237698, -1.0540398, -0.1392331, -0.5084452, 0.5201884, 1.4256452, 1.6968222, -1.8622437, 2.2606048, -0.4436381, -2.4428632, 2.6185835, 2.5700055, -0.0128000, 1.6298676, 1.9203247, -1.1820877, -1.4730193, -1.4002583, -2.8446276, 0.3069639, -0.9288064, -0.3498036, 1.7190115, 1.5274899, 2.8386028, -0.0113960, -0.2629365, -2.7461224, 0.3584656, 0.5534568, -0.8713228, 2.5718880, 2.3522359, 2.6812452, 2.8997044, -0.3777303, 0.6736234, -0.6703953, 2.1208196, -0.9660507, 1.5472929, -1.1673402, 0.1107814, 0.5038401, 1.2256363, 0.4857326, -1.5108235, 1.7994976, -0.3910948, 1.1667085, 0.9806032, 2.0272130, 1.8164579, -1.0888766, -2.2111701, -1.7491431, 1.5955902, -2.2313944, -1.0001492, -1.7143783, 1.4066700, -1.1402543, 0.6198705, -1.1330799, 2.7740544, 2.0357938, 2.6587831, -0.6324963, -2.0833530, -1.4159586, 2.6656297, 2.9403437, -1.2218230, -1.0274030, 2.1992207, -2.9187851, 2.4413647, 1.0666594, -2.8370514, 2.8491168, 2.3676854, 2.1046013, -2.0265936, 0.0042257, -2.7258986, 1.7138953, -1.4909315, 1.6338181, 2.4415902, 1.6521643, 1.8119628, -0.5905237, 1.6884811, -0.9320134, -0.0296216, -2.2585671, -1.5904580, -1.7446942, -0.4071260, 0.8421532, -1.9225698, 2.8903732, 2.0420525, 2.0070963, 1.4543962, -1.3637048, 1.4631338, 2.1416760, -2.0652501, 1.7956457, -2.4121325, 0.7053391, 0.9611561, -0.1251190, -0.9582916, -1.3633590, -0.5851351, -0.8802685, 0.3390205, -2.6530833, 1.0016986, -2.5857963, -1.8813715, -2.3319534, -0.2722318, 1.8565369, 0.6601836, -0.4454128, 0.1635327, -0.3460957, 0.4999581, 1.1758460, 2.1168039, 1.2119603, 1.8108314, 2.0574427, 0.8166895, -1.2670572, 0.8134933, 0.8260508, 0.2756875, 2.9633423, -2.4901166, 0.9315618, 0.7478924, 0.1480391, 2.6038905, 1.6003340, 1.6895059, 0.0030438, 0.0136227, -2.9256936, 1.2370696, -1.7313851, -0.5996957, -1.3948511, -0.1858462, 0.2172290, -0.4980115, 2.6495789, -2.5218263, 2.1387448, -2.2564097, -0.4852043, -0.5178665, -2.4897932, -1.7847908, 0.5059449, -1.1460036, -1.0672936, 2.7475206, -1.5393412, -2.0078081, 0.1651175, -1.0553559, -1.2780558, 0.6573358, 1.6433007, 0.4490870, -0.7909457, -1.0674894, 0.0449661, 1.2898386, 0.7634405, -2.2031650, 2.7505986, 2.7941328, -2.2300760, 1.4734595, 2.7530482, -1.8931402, -1.9344135, -2.6639866, 0.3662690, -0.3902994, -2.1103234, -1.3793964, 1.6347249, -0.4649262, 2.1240989, 0.3460635, -2.1114473, -2.4642838, 1.9593393, -2.9179484, 2.3946592, -1.5183409, -1.5302172, -2.3990353, 0.2756504, 1.6917792, 2.4689127, -1.7592320, 0.7343748, 1.3867088, 1.6367143, -0.0861609, 2.4654443, -0.6677485, 2.6864986, -0.1956412, 0.5039478, 0.3609448, -0.1753442, 2.0399519, -0.1421409, -2.8211013, 1.1378566, -1.4482169, -2.2358710, -1.1534050, 2.8427236, -0.5222450, -1.3316664, -0.6173622, 0.3171313, -0.0063761, 0.2852331, 0.8019916, 1.4812914, -0.1619449, -0.0948908, 0.7242380, -2.0290425, -1.9576283, 0.1868984, -1.6113081, -1.0023158, 1.1846094, -0.3313942, 0.6209858, -2.9562752, -2.4375759, -1.1357562, -2.9157690, -2.0248169, -1.0877404, 0.8744677, -1.1176234, -0.1565634, -0.3990768, 1.4739629, -0.4946939, 1.9974012, -0.1064542, 2.7350219, 2.2313289, -1.1338367, -0.1582032, -2.1278804, 1.8867603, -0.2617088, -1.9577218, -2.1976235, 1.2540755, -2.8945340, 2.9131673, -1.3835834, 0.4650400, -2.9448293, -1.7128607, 2.6958540, 1.1074889, 1.0810150, -2.4251259, -1.5406262, 0.8194569, 1.3231013, 1.2508464, 1.3931134, -2.9005198, -1.8927749, -1.1488363, -2.4506055, 1.4911155, 0.5146038, -2.9743037, 1.8875133, -1.7534793, 2.2560809, -1.3463427, -0.2073602, -0.8317994, 2.3514660, 0.3440772, -2.0187778, 0.2463541, 1.5467902, -1.9318996, 1.8433417, 0.1209071, 0.7154856, 0.3518136, -0.5927536, 0.2969707, 2.9202521, 1.7895315, 0.6965912, -1.8265275, 2.9822898, -1.4136465, 1.4808098, -1.5452035, -2.6845954, 0.6931445, -2.6556369, -2.8729647, -0.3357207, 2.0480530, 1.6047277, 0.8165175, -2.4229813, -2.3135845, 2.8547945, -0.5238284, 0.4151802, 1.2727284, -1.7484246, -0.7990977, 1.0534492, -2.4400265, -0.3952409, -2.7759362, -1.0209445, -0.0288872, -0.6840933, -0.1507097, 1.7971571, 2.5287698, 2.5416080, -2.1134565, 0.1993146, 1.8136593, -1.6138450, 1.1683200, -2.3712424, 1.7130445, -1.3953789, -0.8815550, -1.7705589, -2.5090357, 2.9782104, 2.1646965, -0.3346431, 2.8023221, 2.2460400, 0.0030722, -2.3788475, 0.3926551, 1.9017379, 2.3478879, -0.3893682, 1.7186940, -0.8113922, 0.1951655, -2.2223145, 1.9311597, 0.1455236, -0.9734578, -0.6569061, 0.1597580, -0.1573591, 0.0115065, -1.8407484, 0.2002664, 1.1821880, 1.1265602, -0.9480664, 2.5740069, 0.7241792, -0.8052767, 2.9107285, 1.9038022, -0.3752289, 1.7059393, 1.6971855, 0.8255818, -0.6152702, 0.6704319, 0.9209096, -0.6014537, 1.6873717, 1.8958240, 1.7890963, 2.7786521, 0.9047730, -2.6025683, -2.8801223, -1.6749036, 0.6889167, -2.7715067, 0.2620781, 1.3286453, -1.4029479, -0.5283498, -2.6757684, 2.0715577, -0.8312968, -0.1615663, 0.2942878, -2.2152813, -0.3032704, 1.5871259, -2.2568473, 2.4769331, -2.6545324, 1.8687332, -1.8052122, 2.9830676, 0.7153752, 2.0871695, -1.9408647, -0.9418767, 1.6130836, -0.4410585, -2.9523304, 2.7495910, -2.4029200, -0.7360571, -2.3414562, 2.9696261, 1.8456427, 0.0401753, 1.1063783, -0.9245849, 0.1777231, 1.5095229, 0.7946806, 2.5929457, -2.0208626, 1.1510018, -2.0196365, -1.2775939, -2.1906746, 0.8308692, -2.4604057, 1.5595467, 1.2394062, -0.7459610, -0.7832497, -0.7177040, 1.7997683, -0.7944898, -2.1960552, -2.3612720, 1.6081694, -1.1260275, 1.4326294, 1.4097964, 1.3483476, 2.9693892, 0.3845247, -1.3031914, -1.8568890, -2.0614373, 1.2740661, 1.3632707, -0.3006799, -0.8564998, -0.5414302, 0.2829597, 2.8123117, -1.6946682, -1.6461472, 0.9138544, 1.9530462, -2.8965908, 0.7729008, -0.3547014, 1.2398019, 1.6975552, 0.3529167, -0.9572409, 1.9410631, -1.9641643, 2.5669352, 1.7933536, 1.6939172, 2.8542863, 2.5572460, -2.9618283, 0.5791518, 1.6763101, -0.5215384, 2.0581574, 1.9315493, 1.6046075, 2.7902567, 2.0397379, -0.4392824, 2.9398937, -1.7976201, 2.9377507, 0.7176958, 2.8212405, -2.8251881, 1.4618571, -0.7368080, -1.3449261, -0.2520162, 1.6102782, -1.0186072, 2.3504526, -0.8341879, -2.7085114, 2.8393387, 1.5673051, -0.9116324, 2.2187634, 2.6995113, 1.6715040, 0.0715665, -0.1117585, -0.7419008, 2.8424601, -1.6209094, 0.5168540, 0.6950143, -1.7410410, -2.2835965, -2.5366803, -1.2861571, -1.1326804, 2.4513919, -2.7536555, -0.1823005, -2.7337988, -0.6164735, 0.4210643, 0.4203676, 2.4978346, 0.6327673, 1.7864299, -1.5173807, -0.3027734, -0.7322909, -1.1004678, -0.7693074, -2.1831571, 2.0938194, -1.8443551, -2.9222616, -1.4954537, -1.0306509, 0.6662168, -2.7048793, -0.8849601, 1.8845195, 1.9965495, 1.5792814, 2.7860449, 0.2961915, -2.0355724, 0.9757099, 1.8712083, 0.5710622, -2.4604761, 0.1724544, -0.6362483, -1.6191875, 0.8653062, 2.3452222, 2.0856001, 1.7331335, -2.0834827, 1.5726415, -2.1745193, -0.5949799, 0.6584317, 1.6597823, -0.9680149, 2.6865636, -0.2072373, 0.6763476, -0.0895641, -1.4009838, 1.8708649, -2.5450049, 1.4253667, -1.0795892, -0.4128711, -2.4195640, 0.0880532, 0.5075386, 1.8717734, -0.5012596, -2.0167402, 1.4247252, -0.3297001, 0.2429445, -0.4399617, 1.7582393, 0.4624781, -1.4553348, -1.7431217, -0.4790066, -2.4664939, 0.8007209, -0.7498305, 0.5852434, 2.4746199, 2.8700996, -1.6778632, -1.7592558, 1.6991923, 0.1720498, -0.4668942, -0.7660503, -0.0319059, 2.0899640, -2.2481089, 0.9199056, -2.4404531, 2.6463164, 0.6288098, 2.1995302, -0.9196432, -1.2369157, 0.4010581, 1.0775010, 0.9716444, 1.7313930, 2.1056163, -1.3653794, 2.3976035, 0.8642974, 1.6997439, 1.0006358, 1.7472152, 0.2129733, -2.3584937, -0.8605210, -1.7775969, 2.6760781, -0.7282644, 1.7892591, 1.9986478, 0.1615460, 2.6413778, -2.2842770, -0.3595186, -1.3054586, 0.3250890, -2.7526372, -0.7118861, 1.7316730, 1.7840134, 0.0437112, 2.2487212, -1.5734240, 1.7101472, -0.3122523, -1.8243753, -0.3861124, 0.1088005, -0.9681068, 2.8488258, -0.5303279, 1.5112807, 2.6983920, 2.9481389, -2.4257752, -0.4030277, -1.7318153, -2.6871256, 1.6960686, 0.0587317, -0.4828656, -1.6426440, -1.2763489, -2.6137962, -0.1122327, -2.0386807, -1.3225292, 1.8480596, 1.7261568, -1.8980361, -1.1526649, -2.3243969, 0.2010109, 1.1829788, -0.9939518, -1.1308677, -2.5683320, 0.4984835, -2.0745876, 1.1421710, 0.3335048, 0.2174756, 2.3895793, -2.1445680, 0.6877277, -0.2579619, -0.6470233, 0.3277633, 0.1629567, -1.2902810, -2.1001846, 2.5430634, 2.5791998, -1.6622846, -1.0092665, 1.2515834, -2.9380841, -1.1289069, 1.2973996, 1.8009796, 2.1007225, -2.8530650, -1.7492611, -2.7522056, -1.7654788, -2.6749807, -2.0530522, 2.1234750, 1.0346311, -1.0681682, 1.6580491, -1.9280577, 1.8313195, -1.5832814, 0.4659030, 2.7472709, -2.5224968, -1.3807234, 0.5648729, -0.6097918, 0.1683151, 1.6980696, 1.8213527, -0.7834076, -2.8396419, 2.0191830, -2.0354761, -0.1394318, -0.0516432, 0.0873335, -2.5290359, 1.1065402, -1.9057967, 2.0628014, 1.3903442, -2.8154782, -1.6234084, -2.1556108, 1.9505588, 1.9564780, 1.0601737, -0.8497403, -0.8652825, -0.5012295, 1.4360880, -1.0505613, 2.6693791, 2.2327607, -2.1405382, 2.0038988, -1.6602590, -2.8357721, -1.1411136, -2.9564666, 2.6350785, -0.0106469, 2.6373362, -2.3453295, 1.8440799, 2.0753941, 0.9343165, 1.6598055, 2.6286503, -0.0275707, -2.3399163, 1.2954237, -2.4849285, 2.6628551, 0.8809183, 1.2612122, -0.4594785, -0.1627927, 1.9943678, -2.1133872, -1.4520341, 1.9665511, -1.0011472, -1.4980719, -0.3785351, -0.9920089, -2.3932413, -1.6677397, 1.5701162, -2.7011080, 2.1463601, -0.5756921, 2.1002396, 1.8471946, 0.8241912, 0.0497906, 2.7815920, -1.3978995, 1.7898193, 0.1120272, -1.5469171, 0.5229757, 2.9876768, 0.5638933, -1.8745741, -0.9163465, -2.3607298, 1.3286168, -2.6971575, -1.5436289, -2.6088877, 1.9350554, -0.8618352, 1.9427984, 0.8628100, -1.0450601, -2.7146220, -1.3841356, -2.7629331, 1.4806104, -1.7206281, 2.1970755, 0.2256459, -2.2026964, 1.5328169, 2.3397452, -1.5655530, -2.8057698, 0.9333270, -1.0006318, -1.5122073, -1.4576024, -0.3133668, 2.1828715, 1.2864538, -0.5467176, -0.3274084, -2.9955105, 1.2872337, 2.4868899, 2.0638640, 1.2567012, 0.9959296, -0.4590056, 1.3280835, -1.9032369, -1.8495415, -1.7334590, 2.4500797, 0.6362550, 1.7466336, 2.7437412, 0.6950279, -1.8308012, 0.3796667, -2.7893669, 1.1528114, -0.2593086, 2.7895398, 0.7581800, 2.3205595, 1.3831634, -1.3004919, -2.0118904, 2.4536195, -1.5086091, 0.7092584, -0.5255278, -1.5565826, 0.7757840, -1.1017942, -0.5580204, 2.4431963, 1.4117809, 0.7547940, -2.4873274, -2.9009331, 2.1931527, 1.5315391, -1.4657168, -0.2008619, -2.2125030, -1.5099691, 0.1907421, 2.8852176, 2.8898009, 0.8400729, 2.6120677, -2.1938432, -1.6985953, -0.4151447, 2.2783547, 2.8020819, -1.8182903, 0.3802345, -1.1113698, -2.6462845, -1.8280799, 0.7871904, -1.0209874, 2.0506174, -1.0770403, -2.9035092, -0.0600751, 0.7803722, -2.8063675, -0.0143795, -1.1238550, 1.3212160, 1.2570723, -2.0925179, -1.7468265, -2.8196591, -0.4606755, 0.9137668, -0.2723353, 1.1745629, 0.0584262, -0.2490869, -1.9074573, -2.8131947, -1.6298034, -2.8848112, -0.9916801, 2.2135936, 0.6687628, -0.9598101, -1.8049825, -2.3151238, 0.5985164, 1.6006524, 1.1536240, -0.6723085, 0.4589331, 0.3422268, 1.6644668, -2.8519268, -1.7186583, -2.0473320, 1.3013201, 1.6436899, -1.7798887, 1.1440170, -1.2456803, 0.9124237, 1.7496909, 0.1405915, 2.5266380, 1.3144594, -2.5995549, -0.1924495, 0.5464680, 2.5540567, -2.5250446, 2.9839403, -1.4038432, -1.1056585, 0.8553864, 0.6138624, -0.2616475, -2.3114510, 1.3726679, 1.3632435, -2.8234783, -2.8441596, 1.2342532, 0.4249851, -1.7423788, -2.0524695, 0.2388397, -2.4288681, -2.6295618, -0.7049517, -2.2876633, 2.3597521, 0.1119688, -0.9516139, 1.8450054, 0.7105349, -2.3299274, 2.0154076, 0.2591050, 2.1214937, 0.2806058, -1.8450187, 0.7682202, -1.9855476, 0.7604997, -0.6935415, -1.5772277, -1.5769540, 0.1078926, 1.6103025, -2.4571953, -2.5523952, -2.6597020, 1.8788907, 0.6332254, -0.7956940, 1.4201843, -1.9159752, 1.9874838, -2.6893321, 0.0989326, -2.7503940, -1.0031824, 1.9080819, -1.6488855, -0.5103512, -2.1059359, -2.4862795, -1.1818505, -0.2124562, 0.4648942, 0.3645358, 2.7919288, -1.8539216, 2.9530683, -1.4227054, 1.7224160, 1.8469495, -0.0415033, 1.0772883, -2.9193105, -1.3339881, -1.7632678, 1.7991593, -0.7113398, 2.5556675, -1.9268177, 1.1664688, -1.8128560, -0.8428539, -2.2776065, 1.0591078, -0.0966245, 0.6290160, -1.2630540, 2.8456983, 2.6187685, -1.0464992, -1.8194711, 2.4098612, 0.1050964, -1.5690787, -0.3199687, 1.2975888, 0.6445642, 1.3467526, -2.3324145, 2.9419267, -1.8666542, 1.9345838, -0.1012886, -0.2758907, -1.5326920, -2.4785940, 2.4145827, 1.3990537, 1.9003500, 1.3286612, 1.7595005, 1.9672782, 2.1057574, -2.6680427, 0.6424351, -1.8092060, 2.8082187, -2.3141232, 2.4996332, 0.8355906, -1.4370142, -2.5042480, -0.3431596, 1.7457295, -1.2542560, 0.2750633, -2.9528392, 2.5680868, -1.4174328, -1.4579360, 0.3938584, 1.4675634, 0.8144023, -2.8485483, -0.5976829, 0.1294759, -0.6353294, -2.2986560, 1.8505166, -0.2865710, 1.7942692, 2.5289349, -1.3310483, -2.3655755, 1.2805245, 2.5281122, -2.5544963, -2.8677627, -2.5012809, 0.3638230, 2.8145037, 1.6967550, -0.8934920, 2.4259124, 2.2171274, -1.3112610, -0.9028057, -2.8546222, 2.5295247, -1.8149310, -1.4101109, 0.2745520, -1.2808498, 2.6680889, 2.3070414, -2.0979904, -0.9735031, -0.4078416, -0.6511198, -0.5675718, 0.1703330, 1.8193717, -2.9293340, -1.9118070, 0.4391082, -1.1535271, 0.5509381, 2.1902295, 0.4940383, -1.2738693, -2.8092100, -2.5172006, 1.8403913, 1.4922154, -1.3215106, 0.3525104, -1.2903197, -0.8892532, 0.9677778, 0.1719924, -0.8863006, 2.4810366, -0.4180415, -0.8425580, -2.2830382, -2.6283609, 2.4004580, 2.5887416, -0.3314919, -2.4109312, -2.9639474, -2.1264869, -1.0180925, 2.2723438, -0.9302325, -1.5941933, -1.4538566, -0.5629437, 1.3958572, 1.1962535, 0.1710288, 0.0697708, -0.8550549, 2.6425969, 1.1796467, 2.6726389, 0.9349137, -0.0858386, -0.0686254, -1.1702590, 0.2546891, 1.8592596, 1.6225552, -1.9284029, -2.0034601, 0.2005447, 2.7963844, -0.3973512, 2.9789639, -0.3575333, -0.9372978, 0.4898706, 2.7721463, -2.7729544, -2.6784238, -0.4423938, -2.1713262, -2.5639309, -1.7565127, -1.3405399, 0.5432520, 1.3705207, 2.7772902, -1.0905258, 0.6598497, 2.8226807, -0.8652976, -0.0232251, -0.3445152, 1.1093274, -2.5398375, 1.3518639, -1.1368564, 0.6023576, -2.1002079, -0.1119189, -2.6875382, -1.1990806, 2.6731461, -2.0722327, 1.4645588, -1.7521919, -0.2790822, 0.9679603, 0.2862345, -2.1772721, 0.0544260, -2.6535536, 2.4237446, -0.5629301, 2.9859668, -2.6014064, 1.0728739, -1.4377269, 0.9241883, 1.2898433, -1.6685538, -0.4234545, 0.6271641, -1.0306896, 2.9684255, -2.0278316, -1.1825403, -2.5061909, -1.7792148, 0.3961207, -2.1023197, -0.2041986, -0.2108193, 0.5980079, 1.6092845, -2.6318785, -2.8993262, 2.4240659, -2.6632366, 2.5022182, 1.6616439, -1.7133606, 1.2916928, 0.3286938, -0.5117920, -0.0628178, 0.6799785, 2.2639413, -1.3729097, 1.4319662, -2.6586133, 0.4809785, -0.1518911, -1.6543513, -0.7712342, -2.9352925, -0.0059647, 0.6547870, 0.9611157, -1.5695246, -1.8441572, -1.5983634, 0.5389939, 2.6391592, -1.5030710, 0.8462378, 0.8177687, 2.3185639, 1.2411857, 2.9460955, -0.6838871, 1.7660250, 2.2484063, -2.7554733, 0.7031077, 0.7547130, -0.3088599, 2.3835401, 0.5262556, -1.7056681, -2.5692603, -0.1206035, -2.9038981, -2.0206450, 1.4593769, -1.9186275, 1.9035023, 2.3739311, 0.0865858, 2.2362012, -2.9059718, -1.1421017, -0.8861069, 2.4448211, -1.5415145, 2.9795920, -1.8074760, 0.0734713, -1.1777977, 1.6414817, 1.3477157, 1.6634925, -1.3550114, 0.4708294, -2.8260130, -1.7459776, -2.6759815, 1.9654451, 1.0897543, 1.9103687, -0.5816483, -2.1044358, 0.5401788, 2.0109144, 0.9249352, 1.1192304, 2.6642209, -0.7295016, -2.5327719, -2.7462086, -2.6403738, 2.5832854, -1.0472828, -2.9310556, 2.8627074, 2.0711517, 0.9890635, 1.7049683, -2.3211934, 0.0612214, 0.1596046, -0.4593898, -1.4729096, 2.0811853, -1.4302606, -1.7327350, 1.8077791, 0.1892175, -1.4408872, -2.6167675, -2.0649145, 2.9183698, -1.5958921, 1.8219147, 0.3616349, 2.2249749, -0.7643954, 0.0768421, 2.4495585, -1.5858457, 2.8931471, 1.3217598, 1.9470572, 0.5482814, 0.9724057, 0.6867506, 2.8239281, -2.5891478, 1.4873745, -2.6291697, -1.6076086, -2.0439095, 0.9581399, -1.9364204, -2.9252549, 1.8198457, 1.6338567, 0.0796495, -0.4620770, 1.3600572, -1.0917868, 2.5799671, -0.4182816, -1.5884382, 2.4275401, -1.6971725, 1.9468321, 1.2342086, -2.4404061, -0.3257267, -1.6675524, 1.7431367, -0.9451302, -1.8721925, -0.2851200, 1.1843549, 0.4454712, 0.3581649, -2.3127821, 2.7801466, 1.1716621, -0.3671308, -1.6428925, -0.8411976, -1.6890051, -0.6412932, -0.9620219, 1.4677520, 2.7242892, 1.3494121, 1.3554371, -0.6770964, -0.2371427, 1.0851759, -1.0108525, -2.1257570, 1.7222653, 0.7310592, -1.7590435, -0.0326005, -2.2841801, 1.6176372, -2.1125477, 1.6099510, -1.4274256, 0.5446239, 1.7950845, -2.6581884, -1.0151960, -1.9550257, -0.7585036, -1.2958172, 1.5812789, 2.6501158, -0.2309795, -0.9198090, -2.7227409, 0.6292592, 1.2490038, -1.3263803, 2.4208884, -0.4893857, -1.2648557, -1.5251671, 2.7444056, 0.9582772, -1.9017197, -0.9101549, 0.9938374, -2.8117798, -2.4414510, -2.6807774, -0.2703063, 0.0493513, 0.7987112, -0.1614623, -1.5605153, 2.5142043, 1.6383018, -2.0979021, 2.6354856, -1.3169655, 2.6710446, 1.0411109, 2.3097915, -2.3449888, 1.7542947, 1.8119751, -2.4677928, -2.3462895, -1.0855897, 1.5665649, 1.1164614, 0.7613127, -2.8577063, -1.7069129, -1.4572789, 0.8924944, -2.7131687, -2.2283727, 2.7830696, -0.5087162, -0.7821831, 0.4845899, 0.2215605, -1.8585986, -1.8467579, 2.5580776, -0.6938654, -0.6003693, 0.5492847, 1.5868859, 2.3822286, 2.3745438, -0.6540726, 0.8262244, 1.7908359, 2.2559454, 2.3854418, 1.1898434, 0.2513710, 0.5488103, 1.5611752, 0.5652236, 2.8608537, 2.8330136, -1.4795796, 1.4472153, -1.9030753, -1.9331016, 2.6661830, 1.8704315, 1.7954672, -0.0504216, -1.9049253, -0.4642990, 2.1675376, -1.3896201, 0.0871199, -0.4901600, 1.3273641, -1.3928078, 2.9216522, 1.9988335, -2.8277579, -1.0729047, -2.3600949, 0.7029902, 0.3721535, -0.2699453, -1.0252861, -0.1440920, 0.0325390, -1.2334260, 0.7926420, -2.9044234, -2.3142067, -1.0773807, -1.3689147, -2.1416510, 0.7851611, 1.2708220, -1.9189438, -0.4317213, 2.9119152, -0.0724287, -1.4380482, -2.2217062, 2.2150057, -0.8036699, 1.0837659, 1.8578987, -0.5717914, -2.6111177, -1.9327906, 2.7403401, -2.1615561, -2.5999636, 1.2593024, 1.6747428, -1.2679277, -0.9814593, 2.4291690, 2.7328278, 1.8545751, 2.9884411, -2.7762165, -2.3427364, -2.3236745, 1.4696406, 2.8103505, 1.0582905, -0.9675728, -2.0111337, -0.5611319, -0.5431038, 1.3528500, -2.0129357, 1.9603926, 2.6361081, 2.4521972, -2.7267706, -1.5639384, -0.4934412, 1.7009696, 0.4583962, -2.8844160, 1.3027228, -1.9694593, -0.0078751, 2.7253591, 0.1802678, -0.4234833, 2.9333426, -2.6734593, -2.8352195, -0.9899919, -2.1801705, 1.7300407, -1.7881221, 0.3821823, -1.5644288, 1.7666439, 1.3113170, 2.8011736, -1.9733873, 1.9063418, -2.3739077, 2.8935323, 1.6522036, 1.5312642, -0.9112359, -1.4549332, 2.5891692, -1.9263548, -1.3214228, -1.1966429, -1.2601861, -2.7922900, -1.5190369, 2.9328535, -1.1892206, -2.7787645, 0.4403933, -2.7294333, -1.6307735, -2.3270288, -0.3114869, 2.7265838, -0.6837065, -1.1581722, -0.3091122, -1.3996502, -1.3736990, -2.0533840, 1.1101445, -2.1821069, 2.7052916, -0.7000091, -1.3765222, -2.5463227, 0.7380282, -2.7760765, -1.7909212, -1.3904857, 0.9586628, 1.7251215, 2.0021335, 0.3383145, 1.6603706, 2.1897762, -0.6374900, 1.3165081, -0.6887095, -2.6080997, 1.5866676, 2.9276726, -0.3368274, 1.3492956, -1.8489167, -2.4839657, -2.8115008, 2.1068299, 2.3497712, -2.6971445, -2.3611929, -1.0920726, -1.4453137, 1.2390879, 1.0702936, -1.3266603, -2.4297820, -1.4492042, -0.3630782, 2.0485853, -0.1425653, -1.9488460, -1.3321093, -0.3392952, 2.4918001, -2.2825380, -2.8968140, 1.8485882, 1.2661319, -2.4204567, -2.9548106, 1.0775582, 2.6227658, 1.5272496, 1.5895058, -1.3802561, -1.1901212, -2.3052029, -0.6077759, -0.0631239, 0.2575414, 2.0158087, -2.8145985, -2.6821468, -1.7861501, -1.9505316, -1.8382903, 2.3418999, 1.3127844, 1.8718363, 2.1702039, -2.4032628, 0.5688814, -1.3102946, 1.1241865, 2.1121315, 1.3484082, -0.6739761, 1.9718761, -1.7608540, 2.1491762, -2.6656516, 2.2046790, -2.8260635, -0.8471858, 0.7270164, -0.3779318, 2.3605430, -1.6964700, 1.5981426, 0.8478840, 1.4844817, 1.7377267, -0.7494685, 1.7171738, -0.8870953, 0.9982999, 1.1764285, 2.6890476, 1.7773676, 1.4225654, 0.3510898, 1.6828686, -2.7912499, 2.3674576, 1.3660439, 0.8132901, 1.1392083, 1.0979124, 0.3760555, 2.9083413, 1.3367980, 1.0028480, 0.2063951, -0.8517681, 0.8892718, 1.2822375, 2.9013282, 0.4942881, -0.5196317, 1.1977092, -2.6923299, -2.8608836, 1.0747173, 2.9283632, -2.5993128, 0.9339501, -1.7287551, 0.5888916, 2.9646050, 0.8451709, 2.8633771, -0.1449145, 1.2925603, 0.2868373, 1.5038944, -1.3474672, 0.0639273, 2.3519689, 1.4519224, 2.2625754, 0.6959814, 0.4980636, -1.6478718, 2.6480578, 1.9778886, 1.4300914, 2.4587738, -1.9256438, 0.7380295, -2.9790918, 2.0160562, -0.4680390, -1.7640535, -0.4281436, 0.1683705, -1.3991584, 1.1001124, 1.1613241, 1.4782974, -2.2584376, -1.9990369, -1.6953720, 2.9947415, 1.1471421, 1.5346807, 1.4815676, -2.3331198, -1.6868205, -0.7782222, -0.8775254, 1.2577051, 1.8468279, 2.0035833, -0.8977331, 1.8414745, -0.5341238, -1.5015796, -0.2705174, -0.3672537, -0.1218927, 2.6980535, -2.6285580, 0.1700808, -0.1671113, 2.9884021, 1.1530660, 0.7484201, 1.1638787, 0.6210520, 2.7269914, 2.3449113, -2.7252646, -0.6611947, 0.1277309, 2.4340692, 0.8723924, -0.9663505, 2.7207868, -1.1665049, -2.9691658, -2.7167822, 2.9530431, -0.6599550, -0.9934385, -1.7871552, 2.2190969, 2.9584299, -1.8336236, 2.4517922, 2.2364391, -1.7727013, -2.4236212, 1.7668605, 0.3107494, -2.1137754, -2.3649082, 2.7435891, 2.0155078, -2.3442745, 0.0990466, 1.0320955, -2.7736892, -1.5140921, 2.2440537, 0.1615298, 0.7084499, 2.2497816, -2.1277081, -1.6048340, 2.4333250, -1.2041911, 1.1484027, -0.1621639, 2.2666271, 1.9922068, -2.3001991, -0.8005702, 2.8444784, -0.7069769, 1.5102222, 2.5198682, 2.3008850, 2.1972851, -1.9622990, -2.9613469, 2.0694491, -0.2284345, 2.7847851, 2.3011260, -2.1279632, 1.8073920, -0.4372860, -2.1006063, -1.3668369, -0.6554556, 0.9486633, -2.3566530, -1.8663441, -1.8991499, 1.2008044, 2.6183408, -0.0660482, 2.3218413, -2.7064522, 2.9949808, 2.8163085, -1.3944855, -1.8318213, -2.9815813, -0.2446423, -0.8117706, -0.1054793, -2.4968435, 1.2566538, -0.5353004, 1.6207372, -2.4167499, -1.1987452, -1.1725075, 2.8590855, 0.7860423, -2.9382027, -1.7198495, -0.3549850, 1.4549472, -0.9166502, 1.2406085, 2.9785137, 0.7493751, 0.9762897, 0.0319879, 2.1785631, 0.8305303, -2.4078969, -0.4557930, 1.6981611, -1.5416001, -2.5316798, -2.2090114, -2.3622461, 1.7271179, -1.3149357, 0.5640522, -0.5615485, 0.3602706, -1.7539399, -2.2138771, -0.2634426, 1.9468947, -2.4006654, 0.9803912, -2.6693433, 1.4249481, -1.0191825, -0.8417840, 0.0797557, 1.8357629, 1.6920700, 0.3237870, 1.7653981, 1.3987066, -2.4403729, 2.8229761, -0.3455639, -0.3438170, -1.2308389, -0.2361643, 0.6616311, 1.9537282, -0.9404842, -1.8032403, 1.4385446, 0.0832129, -1.9154519, 0.2101012, -0.0591138, -0.8558929, -0.5420487, 0.6147347, -1.3501550, 0.9223968, -1.4893551, -2.8274039, -1.7384289, 0.4739164, -2.7850073, 1.6860029, -2.4289962, -0.5772748, 0.7569370, -0.0123966, -1.7272255, -1.4017637, 2.4084478, -0.7608691, -0.3865078, -2.5486106, 2.8795454, -0.0819213, 0.3668178, 2.8946718, -1.8567458, -0.5078529, -1.5493102, 2.6143112, 2.9473705, 1.5957247, 2.3356732, -2.1592234, 2.0869672, -0.1238974, 0.1716869, 1.4342805, 1.6882020, 0.7515862, -0.0415504, 2.5197992, -1.2321700, 0.3354297, -2.4015741, 0.9763453, -1.8702584, -2.6363325, 0.4981670, -1.6361197, -2.9320863, -2.7896906, -0.7278110, -1.7178120, 2.5279390, 1.7587909, -1.9492449, 0.8045875, -0.4285579, -1.8744214, 0.9485483, -0.0384506, 1.4420274, -0.5428229, -0.8847680, 0.8523779, -1.2633963, -1.0020008, -1.6072980, -1.7466671, 0.6198824, -0.0304512, 0.8192925, -2.6060462, 2.4764959, 1.0008964, -2.1655564, 2.4827676, -1.9939723, -0.4868492, -2.6409309, 1.2275578, 0.7860667, -0.3749009, -0.1296546, -2.0169705, 2.3179198, -2.7789960, 2.7281364, -1.6306209, 1.4278892, -2.4193438, -2.0813327, 0.8115133, 1.2798094, -0.0742169, 2.1705114, 2.7164953, 0.9821761, -1.0476125, 0.2619420, 1.0812024, 2.0716657, -1.3412075, -1.1248821, -1.6686746, -0.5001357, -1.1506616, 0.3500098, -2.6901652, -1.0866440, 0.8712451, -1.8212883, 2.5317308, -1.9260054, 0.5270882, -0.9377332, -0.4513217, -2.0463387, -0.6984431, -2.1272549, -0.6006678, 1.3586869, 1.4834113, -0.3323088, -1.4668735, -1.0972776, 2.3745271, -1.1283578, 0.8874077, -1.0377692, 1.1023773, -0.7856243, -2.9153846, -1.5338009, -2.6230134, 1.9726493, 2.3794258, -1.8351788, 2.4429975, 1.5907245, 1.1066277, 0.9206081, 2.9413887, -2.3129333, 2.9883565, 1.4720237, 1.5757420, -2.0936126, 0.9267466, -2.0290705, 1.5442827, -2.4351367, -2.8714140, 1.2069352, 2.9914421, -2.9141648, 2.8732751, 2.4804046, -1.0767993, -2.7913549, -2.2220982, 0.2911926, 2.1732417, -2.9660743, -0.3903164, 2.1171929, 0.0367984, 0.3529198, 0.8092620, -2.7549213, 0.6984564, -0.4739676, 1.7302002, -2.6126420, 1.4445762, -1.8897992, -1.2538841, -1.6952229, 1.7019172, -0.6383084, -2.6244204, 1.2797415, -2.1482788, -2.4655842, 2.5196004, 2.7775283, 2.0480636, -0.5739715, 2.2895690, 0.9703181, -1.7824419, -2.4672935, -2.1568162, -0.3288941, -0.4254316, 2.2986748, 2.8718351, -2.8703927, -1.8604186, 2.5238960, 1.3261251, 2.1951198, 2.1083291, 2.0132511, -2.5979804, -2.2612142, 0.8431135, 2.0713938, -2.8380785, -0.8572747, 2.3119020, -1.8319865, 2.8997962, -0.6388207, 0.1161874, -2.0330492, 1.6199985, -0.0949730, 1.8298233, -0.4120283, -0.7167007, -2.6472053, -2.6101354, 2.6754702, 1.5644574, 0.9380472, 2.7506345, -2.8946102, -1.9004825, 1.9407012, 0.6572658, 0.9289347, 0.5503878, 1.8333177, -2.1987308, -0.4451889, -1.7147021, -0.3654777, 0.9934452, -1.9224433, 1.6186925, 0.7239059, -0.5199707, 2.2432001, -0.0849249, -2.2245515, -1.5114703, -2.0791073, -2.0321009, -0.7441795, 0.1891809, 0.5865817, -0.6857163, 2.3004784, -2.6790240, -2.0305691, 1.9405177, -2.9064349, -2.1268057, -0.5421224, -2.1398140, -2.0132682, -1.3690306, -2.5334822, -1.9403980, -2.7686538, -1.9081114, 1.8835772, -1.8170066, 1.2070035, -1.6243106, 2.3528132, -1.1268382, 2.4640522, 2.4841035, -2.6184836, 1.8662640, 2.1120676, 1.4380724, -0.2130874, -1.3894509, 0.1161460, -2.5414006, 1.8613039, -2.9587559, -2.8398847, -2.7729833, -2.2305103, -0.1388146, 1.0078638, 2.7870456, -1.4036156, 0.9449841, -1.3245553, -2.9312179, 0.0075762, -1.7650034, 1.5270464, 0.3438461, 1.5325916, 1.5496091, -0.0676711, -0.3590711, 0.3629450, 2.2944874, 0.0246575, 2.7375404, 1.7617361, -0.1842502, -1.4591982, 0.7841828, 2.6286611, -2.5369215, -2.7801929, 0.5259904, -1.7738906, -0.0255729, -1.0558421, 1.8919582, -0.5460403, 0.0036820, -1.0157450, -0.6263910, -1.9024330, -1.6767118, -0.9866393, -1.1432124, 2.7042909, -2.2696345, 1.3393138, 0.9618892, -1.2585371, -1.3986117, -1.3809043, 2.2435855, 1.0274099, -2.6002470, 1.6020275, -1.2419733, 0.8318456, -2.3792662, -2.9594257, -2.3726974, -1.6037455, -0.6364196, -0.1729657, -2.4532788, -2.4555521, 1.5916838, -1.1421578, -0.2166940, -1.7085402, 0.1744559, -0.3385207, -1.1390236, 1.6998429, -2.3520052, 2.0408126, 2.8445393, -1.5028674, 1.6711801, -1.7349976, 2.9421887, -0.2961188, -1.5434508, 0.3466087, -1.4039157, -1.9780102, 2.6291500, 0.7543686, 2.6521655, -2.9838860, -0.9486500, -2.7191948, -2.9684628, 0.7562189, -1.5447516, 1.5435225, -0.2598304, -2.5656140, 2.6503287, -2.7938810, -0.1019416, -2.3866557, 2.9563606, -1.3734051, -1.8910962, 0.3282254, -0.7452423, 0.5361603, 1.7187268, 1.0471317, 1.9506403, 2.4870903, 2.8992515, -0.8298513, -0.2503045, 0.4466889, 0.7833319, 1.8210880, 0.9176625, -2.3861008, 1.9885665, 1.6825365, 0.4278681, -0.0379228, -0.7899916, 1.1696621, -2.5402250, -1.5129573, 2.3431520, -1.7440498, 0.0115363, 1.4677982, -2.2083455, 2.0304556, 0.4777263, -2.3119058, -1.8871962, -0.0010890, -1.2612695, -2.9284864, -1.2997670, 2.1828070, 0.2585156, -1.2632303, 1.3963281, -0.8790856, -1.0355326, 1.0237856, -2.3287068, -2.3093713, 2.6516827, 1.3147695, -0.3627111, -1.3076243, -2.8841109, 0.6676982, -1.9931050, 0.2153270, 0.5046263, 2.8686477, -2.4363660, 0.1853894, 1.5516079, 1.5464594, -1.5660134, -0.9524094, -1.9812567, -2.3611290, 1.9471348, 0.9507919, -2.9138502, 0.5587991, -1.3042014, -2.9745453, 0.5280521, 1.7717592, -1.3902000, 2.5029298, -1.1664632, 0.9579095, -2.4233330, -0.5648300, -2.9944147, 0.3238568, -0.9339407, -2.1878382, -2.5869956, 1.1902586, 0.8981368, -1.1552665, -2.1402682, 2.5728062, -0.8079380, -2.4477329, 0.3682016, -2.8860306, -2.0529517, 0.6608439, -0.8800991, 1.9766687, -0.8750849, 2.0512725, -2.9282494, 2.3647703, 2.2255859, 2.6563527, 2.0266608, 1.4812354, 2.4429693, -1.5730151, 0.1009874, -0.3324976, -1.3527255, 2.2057585, -0.2999150, 1.2235450, -2.1257678, 0.2651106, 0.5622272, -0.6535911, 2.3271016, -2.5590821, -1.9846908, -1.9870448, 1.4267418, 0.8859607, 1.2415230, 2.7312581, -2.2670406, -2.8849659, 2.4130110, -2.3929549, -2.9878847, 1.1619957, -1.2100777, -2.2940264, 1.9812340, -1.2026626, -2.7251366, -2.1327389, -1.2179615, -0.0989886, 1.1109581, -1.6978504, 2.0824377, -2.7373792, -1.1394664, -2.6060101, -0.6660345, -2.5627164, 2.9762771, 2.9712346, 1.2696589, -1.4724055, 2.8071556, 1.2321561, -1.6541081, 0.3668601, -2.0326364, -2.8943078, 1.9554738, 0.2936098, -0.6675709, -2.1911529, -0.0015894, 2.0561056, -0.9435450, -2.7646773, -2.2982471, 1.2155834, 2.6229186, 1.2278240, -2.0059110, -1.6635109, -2.5977971, 1.7968091, -2.0082246, 2.4727232, -0.0825464, 2.2002569, -2.1737758, 1.2366287, 1.2473665, -2.0667973, 1.9544017, -0.8071553, 0.3833252, -0.9397746, 1.7701130, -2.6631551, -2.1819630, 1.2511123, -2.4425745, -2.5985558, -0.6932676, 0.3746705, 1.4744281, 0.2516712, 2.2865572, 1.3785425, -1.1388536, -0.6673346, 1.4982465, 0.2228458, 1.9617619, 0.3618248, -1.9154532, 1.2028193, -2.3701840, 0.5416955, 0.7631094, -2.3174248, 0.7162890, -1.1669554, 2.0819767, 2.9685634, 2.8399942, 0.5437160, -0.7825133, 1.1054414, 0.4115190, -0.3366731, 2.0555443, -2.5455470, 0.6465669, -0.1766795, -2.4913877, 2.3555044, 1.8685724, -1.6857954, -2.7055060, 1.7003035, 0.9309468, -2.1300776, -1.9075295, -0.2645610, 1.7393988, -0.7045317, -1.8352123, -0.5051571, -2.9737206, -1.5427700, -1.7528988, -2.6185858, -1.1374149, -2.1077075, 0.5012312, -2.8889589, 2.6476285, 0.7106937, 0.3259722, 0.6745765, -2.4606141, -1.3883440, 0.6302868, 0.1923986, 1.3172777, -1.9973868, 0.9806589, -0.5765862, 1.4067251, 1.9898538, -0.9315710, 0.1996032, 0.2276020, -0.3957851, -1.8139992, 1.6298489, 1.2811700, -1.5099262, 1.7145623, -1.1209761, 2.4790935, 0.6297366, 0.2259282, -1.2600729, 0.0361781, -1.3249709, 2.7172158, -1.2469560, 1.6363849, 2.8169918, -1.3676415, 0.3630195, -0.0051645, 2.3551340, -1.9543944, 1.0227825, -1.5570316, -0.7347793, -1.9473042, -0.8425916, 1.3935935, -1.5225851, -1.5937846, -2.9836614, 1.9567696, -2.7509344, 2.2265047, 1.4424435, 1.6291811, -2.2476795, 0.9017014, 2.9836188, 1.2977387, 1.9299492, -0.9659448, -2.0510199, -1.3870825, 2.6638430, -0.2803667, -0.1919282, -1.1623952, -0.0145528, -0.8808717, 0.8208253, -0.4247849, 2.7037288, 2.4514688, -1.5336502, -0.4002591, -2.3633623, 2.6006016, 2.1617131, 2.6796831, 2.7995314, -1.1462005, -2.2725653, -0.5686007, 1.0139096, -1.3722720, 0.7623249, -2.4151569, -2.4602166, -2.8595730, 1.0958787, -2.1366250, 0.8929888, -2.5300946, 2.4232203, 1.5799590, 2.1441114, -2.2724999, 1.8910269, 0.1611220, -0.4233376, -1.1848431, -2.8009223, -1.8741394, 1.9021103, 1.2422332, -0.9312547, 1.8969849, 1.6386492, 2.4705258, 1.0167276, -1.8450494, -1.8654637, -1.1368821, 1.1571465, -2.9875167, 2.0266903, -0.4623640, -0.4272305, -1.5042440, 0.6063296, 1.1674599, 1.6736737, 0.6686448, 2.8823109, -2.3675217, -2.3805527, -2.6099698, 0.5405538, -1.5017103, -0.0838816, 2.7900711, -1.4769376, 0.2488520, -2.6618342, 1.8815910, -2.6828563, -1.6386973, 2.1559443, 1.6248710, -2.7373947, -1.3566790, -2.7610465, 0.7892861, 1.5611345, -2.1767946, -1.0582533, -1.5779425, 1.3461663, 0.7538014, 2.2479511, -2.0495012, 1.7481719, -1.4971591, 1.3782792, -1.9064582, -1.5584943, -2.7672980, 1.2347545, 2.0951162, -2.9014490, 2.6806087, 0.1733654, -2.4897732, 2.5711322, 0.4175564, -2.2084433, 0.1058869, -2.9252667, 1.6499860, 2.6812068, -2.7067659, 2.6668399, 2.7624073, 0.8117463, 1.9128900, -1.8445686, -0.9497904, 2.1079938, 0.9112661, -0.1744071, 1.7146323, 2.1840238, -1.8195612, 2.2776993, 0.2690840, -2.5425187, 2.3500821, 0.4285043, -0.9208464, 1.4925366, -0.8088606, 1.2623470, 2.8079298, -0.3100017, -1.1273747, 0.8982299, -0.6459093, -0.4214128, 1.8674959, -0.7231923, 2.4138453, -2.6305340, 0.8235889, 0.5240426, -1.6322456, 1.8085997, -1.2028314, -2.1989098, -0.0696857, -0.3998124, -2.6421542, 1.5298886, -0.4837358, -0.3195471, -2.7335659, -0.9408162, -0.7576195, -0.7793926, -2.8169459, -2.7186081, 2.4911349, -2.9021211, 1.9744261, -1.6903146, -2.0645422, 1.5622661, 1.5331922, 2.6690329, -2.1394074, 0.9684678, -2.3492579, -0.3443362, -1.0622788, -2.0889796, 1.6686463, -1.3542708, -1.7577165, 0.7066097, -0.7995878, 0.1424235, 2.0380672, -2.3349948, 1.9937117, -0.7619616, -0.4512729, -2.7778030, 1.3582643, -1.1490500, 2.7011330, 0.9267385, 1.5426027, -2.5958384, 0.8304446, 1.3008654, -0.9500038, -2.4780378, -1.6370039, -1.1840819, 0.6603069, 2.1573290, 1.1419812, 0.6581926, -0.3304953, 1.4630208, 2.4939038, -0.2635497, -1.1090863, 0.9722327, -1.6000767, -1.8312265, 1.3229132, -2.9398476, 2.5113901, -2.1892518, 2.2056257, -0.9956345, -2.1925464, -0.7902831, -0.8225819, 1.1426060, -2.9123519, -1.8483490, -2.4804188, 2.0673176, -1.0247913, 2.3530386, -1.6137618, -1.9950068, -2.0993338, 0.0552678, -0.3810327, 0.9408055, -1.2163529, -2.2820735, 2.2278501, 0.7958507, -2.9274894, 0.3808746, -2.1096913, 2.9650209, 0.3936367, -1.4112822, 2.8653554, 1.6136892, -1.8045746, -2.8106536, 1.9164664, -2.5865967, -0.4999737, 0.3171732, 0.6083496, -0.9319726, -0.8676233, -0.4519955, 1.5722917, -2.0625833, 1.1442406, -0.6813315, 0.5401216, 2.2726209, 1.0692296, -1.2490312, -0.2021682, -0.9384290, 0.6066031, -0.9091391, 1.8969384, 0.6991653, -0.9155247, 0.8762903, -1.3094872, -1.8456772, 2.1714530, 0.9280887, 1.2969145, 2.0148618, 2.8130851, 1.3174793, 1.6598023, 1.8460587, -2.3881120, -1.0503940, 0.2791169, 2.9678186, -1.9995199, 0.6423192, 1.4742872, 1.7006967, 0.1278898, -2.2751395, 0.0771037, -2.1938354, -1.3029326, -1.1328501, 0.9741827, -0.9970554, 0.2124192, -2.3930018, -2.4422341, 0.5154326, -0.1694175, -0.9095934, -2.3531616, -2.8162759, 0.5476245, 1.2695957, -0.1299749, -1.3635239, -2.2887186, 1.2253011, 0.1646931, -1.8718846, 1.6011329, -2.4479980, 1.4662741, 1.8646666, -1.5955451, -2.6751613, -0.2652444, -0.8625089, 1.7813197, -1.8303455, 2.6714539, -1.2812467, 2.4357448, -1.3808501, 1.4313005, 2.7471452, 1.2269339, 2.7765494, -1.0985854, -2.7308180, 2.3802374, 1.2030964, -1.6666636, -0.3018421, 1.2083491, 1.6578844, 2.8940005, -1.9362598, -2.1566677, 1.3423947, 1.2626704, -2.0634417, 1.0460535, 1.2333422, 0.8296633, -1.6163465, 1.8534852, -0.1890203, 0.0850697, 0.3689421, 0.5569142, -0.9311866, 2.9826888, -2.3674340, -2.6980708, 1.6383044, 2.2783560, -1.7283067, -1.0240949, 1.7390725, -1.5115630, 2.7357136, -2.2175839, -2.7349331, 1.9014680, 1.4020523, 1.7781018, -1.2477516, 1.2966555, -1.8655089, -0.0197456, -2.2206906, -1.0771008, 0.1430785, 1.9031360, -2.8836477, 1.7628989, 1.3738674, 2.2356824, -2.7648235, 1.7644940, 0.8496512, 0.4728743, 1.8823197, 0.6846036, -1.3314738, -0.6938388, -2.6592035, -0.0858265, 1.9579846, -0.2130055, -0.6202324, -1.3542341, 1.3811203, -2.9807734, -2.3953697, -0.3731196, 1.8158289, -2.9041405, 2.6918733, -0.4027897, -2.4287255, 1.1937236, -0.8184809, 1.2997253, -1.0976764, -2.4940791, 2.1130785, 2.4177183, 1.1438334, -0.2593352, 1.8231234, 1.8334061, -2.5588950, -0.9683940, -1.8583988, 0.4188210, -1.9190370, -2.8743091, -0.4241935, -2.4414836, -2.5759964, -1.4216368, -2.1527710, -2.5532543, -0.8336048, 1.1271175, -2.6665436, -2.2325040, -1.8337361, 0.2211667, 0.4061846, -2.5505631, 0.9833260, -1.7194049, 0.1750473, -2.8870046, 0.2835757, 0.1506677, 1.4631888, -0.9591655, 2.5486474, 2.3327520, -1.9654962, -1.0155308, -0.3741604, -1.1545803, -1.8416386, 1.1735528, 2.7433123, -0.2194200, -0.5555242, 1.9974873, -0.5728536, -0.9694558, -1.8391639, -0.3449863, 2.1897574, 2.0052730, 0.1245544, 1.9101056, 0.7450166, 1.7519026, -1.7594752, -2.7146945, 0.8337474, 0.4357039, 1.7331488, -0.5474263, -1.5258753, 2.3025839, -0.2464010, -1.8780044, 0.0975037, 0.1392195, 1.1428693, -2.0483220, 1.5284286, -1.7262780, -2.6403534, 2.1042440, -2.0475188, -1.7721571, 2.4981130, -1.3329879, -0.5153069, 0.2942097, 1.6710626, 1.6852713, -2.5233706, -0.8733278, 1.5116113, -0.5623664, -1.3835155, 2.6339761, 1.9074711, 2.1011038, 0.2421051, 1.9816505, 0.2092778, -2.5722740, 0.9968502, 1.7507763, 2.3783482, 0.4382059, -2.5698040, 0.2820581, 0.4650231, 1.6344265, 0.4555126, -1.3061144, -1.6523903, -2.9234439, -2.1993374, 1.5913925, -1.9194353, -0.6657480, -0.0006236, -2.3228521, 2.5920642, -0.5865400, 1.3692545, -1.4254352, 1.9347560, 2.3778819, -2.1492396, -2.7580796, -2.6606139, -0.6245597, 1.3330289, 1.4133573, 1.0821502, 1.9938788, -0.9665034, -2.3221496, -0.8969478, -2.6359716, -1.4914975, 0.2687094, 2.1778865, 2.2169654, -1.0343250, -2.7742712, -2.7727251, -1.4209093, 0.3288056, -0.3182774, 2.7514775, 2.5640560, 2.1313207, -0.8234765, -2.7949411, -1.7593722, 2.7663618, -1.1212245, -0.9454310, 1.0608400, -1.9443171, -1.8612292, -1.1767906, -1.0330790, -0.0831402, -0.0191284, 1.5258150, -1.7642883, 1.2009699, -2.1362717, -2.4215774, -1.4210309, -0.0812663, 1.1621966, 1.5351303, 0.1525042, 2.6079716, 1.5376115, -2.8569395, -1.7802103, -2.4923914, 2.8890252, -2.1423332, -1.5936665, -0.5367043, -0.2046653, -2.1053246, -2.8130598, 1.1582768, -0.9661985, 2.1262751, 1.1171122, 1.8219689, 2.7450700, 0.2721950, -2.1234124, 2.1042300, -0.9365147, 1.3688532, 0.9905363, 1.1229907, 1.1380944, 2.7537365, -0.9063377, -2.9081405, -0.2828704, -1.4121832, -0.2055195, 2.5303381, 2.7060810, -1.2260081, 1.9851320, 1.2788275, 0.5968476, 2.1909867, 0.6304999, -2.4661176, -2.2379470, 1.6007260, 2.3224859, 0.7967066, 0.0662942, 2.6845464, 1.5817640, 0.8222762, 2.6700487, -1.1529879, 1.1886516, 0.7175720, -0.5646981, -0.4372525, 1.8371333, 1.9055563, -1.9006354, 0.2478012, -1.3130250, -1.9141664, -1.1127690, -1.5750500, -0.5225377, -0.2846382, 2.0688386, 1.5074533, -1.0366204, 1.8296974, -1.2797248, 0.2134227, 2.4253635, -1.4769369, -0.2535760, -1.9646079, -2.1650516, -1.3272786, -2.7919733, 0.3253182, -2.3325632, -2.8537223, 0.3169646, 2.0183891, -0.0704584, -1.0284063, 0.8073419, -0.1787342, -2.8512343, -1.1907794, 0.4418222, 0.8643520, -2.2257507, -0.0810850, -2.7264834, 0.5812420, 0.7058815, -0.9673814, -1.7607353, 2.4408045, -0.6450892, 0.6489583, -2.0411515, 0.1391625, -1.7593377, 2.5432501, -2.8789210, 1.6274040, -1.7629092, -1.1972932, 1.2043681, -2.3467235, 1.8758505, 0.1410344, 1.6481681, -0.5083377, 0.1690078, -0.0846596, -2.1191071, 1.2080498, -1.2769202, 2.8225715, -0.4013895, -2.2994126, 1.4063553, -2.1761678, -0.3499507, -2.9316678, 0.3629932, 2.8368465, -0.3754724, -1.7142925, -2.9949306, -1.1614358, 1.5738075, 0.3710213, -2.8262502, -1.9715043, -2.2487365, 2.1897543, 1.6279127, -2.9222571, -0.9279536, -2.0353967, 0.1592050, 2.6724240, -1.4022840, 0.4916160, -0.8611189, 2.8984553, -0.9180453, 2.0506210, 0.3948725, 2.1144186, 2.2111810, -1.1893819, 0.5061738, 2.2106067, 0.3388705, -0.1717327, 2.2047384, 1.5645200, -1.2105350, 0.4649498, 1.7939683, -2.9510640, -0.6792694, 0.6926012, -2.3599462, 2.2282591, -1.6703589, 1.3404545, 1.4572843, -2.4376742, -0.3781808, -0.8889873, -1.9362457, -1.3999098, -1.3395914, -2.5176135, -0.6076558, 0.7643612, 2.4559759, 0.3917122, -1.0953817, -0.6647482, 0.9805680, 1.6570054, -2.8248059, -1.3789835, -0.4400450, -0.4757478, -0.4247859, 0.5612622, 1.6342064, -0.6522062, 1.3964145, -1.5274016, 0.6721083, 2.7445363, -1.8140654, -1.4387024, -2.5788580, -1.9184302, -0.9678768, 1.3049149, 0.7884385, 0.3878863, -2.8183569, 0.1393650, -1.7282638, -0.6856427, 0.0802149, 2.4931552, -0.2326338, -0.0450228, 0.7700640, -1.0892716, 1.5267775, 0.8611683, 2.4628304, 2.0982809, 0.7485468, 0.0722476, -0.1575181, -0.5539633, 2.9421147, -2.9089744, 2.4740195, -1.4008136, -0.8782888, -2.1696874, -0.8116913, 2.3237115, -0.7366374, -1.5470985, -1.0538352, 0.6247892, -0.2674077, 2.6028745, -0.1147919, 0.6333394, 2.2673642, -0.0308621, 2.8554478, 2.4754745, -2.1987516, -2.7523365, -2.9941802, 0.3868281, 0.3116553, 0.3427153, -1.5714572, 1.9147209, -2.0646441, 2.6489534, -2.2157274, -0.8261538, 0.3103437, -1.1964051, -2.6491794, -0.8265619, 2.0467481, -0.4946085, -2.1836191, 2.3758713, -1.3907530, 0.8690626, 2.8307668, -1.3382347, -1.0084033, 1.6404160, 0.3061126, -0.0663475, 0.0114808, 1.9607636, -0.4111631, 2.5752159, -2.9543696, -2.6896260, -0.6919830, -1.7369236, -1.7862453, -1.1834744, -0.3320141, 2.9836826, 2.6207195, -2.0250339, -0.9139157, 0.6054629, -1.9097132, 0.0463554, -0.1607657, 1.4670396, 0.5326752, 1.8814142, 0.2772430, 0.6170605, -0.2361358, 1.6685731, 2.6765082, -0.6531078, 0.7174854, 1.3083225, 0.1028259, -0.9456503, 1.1122340, -2.2832525, -2.4518148, -0.5915649, -2.3050580, 0.3546187, 1.7847337, 0.0672373, 2.5832731, 2.1124309, 0.2900009, -1.9766859, 0.6515858, -0.9326296, -0.0921457, -2.7265205, -1.5012725, 0.4478243, 0.7093528, 1.8920434, -1.1157577, -0.9998966, 2.4176324, -0.2226870, -2.6447907, 1.0796858, -2.2687312, -2.4381050, -1.3906843, 0.6797019, 2.1342009, 0.7113300, 2.6520446, -2.9961561, 1.4857133, -1.2001523, -1.7323530, -1.8364551, 1.5957591, 1.9213763, 1.7452423, -2.1547706, 2.9801745, 0.9225095, 0.6860509, -1.7735535, -2.0169666, 2.9098909, 2.1363788, 2.5965113, -0.7471675, -2.6839265, -1.0453992, 2.9247477, 2.5355880, 2.8292885, 0.1382970, 2.3489779, 2.5471451, 2.6851712, -2.4371702, 0.6491171, 2.2133673, 1.5631505, 1.5856993, -1.2944340, -1.5857784, 1.9657985, -2.8489023, -2.7170201, -2.9471563, 0.4539209, -1.1124701, -2.1065529, 1.1191045, -1.0502327, -0.9486194, 1.4735565, -0.5237196, -0.3172605, 2.8930628, -2.8713464, -0.4183825, 2.5229905, -1.6742797, 1.4636137, 0.9898283, 0.7699836, 2.3798043, -2.3655296, -2.2181401, 0.3898187, 1.1916155, -2.1652599, -0.5921281, -0.5344185, 2.9963366, 1.9277812, -2.4203236, 1.7994924, 1.2729900, -1.5792443, -2.9082927, 2.6057337, 2.3231530, 1.4003982, 2.1332534, -2.5647966, 0.9615313, 1.9152137, -2.0777559, -2.7640728, 1.1102597, 2.2629704, 2.7046549, -0.2216252, 2.7353085, -0.6411990, -2.5806188, -2.7648432, 1.7344494, 0.3025148, -1.9172447, 1.7203609, -1.4619336, -2.9307152, -2.4553432, -2.6372053, -1.0504707, -1.4317091, -2.6472982, 1.8369951, -1.7265288, -0.2531062, -0.7281305, 2.9788037, 0.8251248, -0.9169451, 1.6252571, 0.2801430, -2.4525932, 2.1605800, 1.5893995, -2.9961989, 1.4343000, -0.0035966, 1.5029961, 2.2496894, 2.5422668, -0.5798418, 1.1175231, 0.4294066, -2.9610234, -2.8088311, -0.8078020, -1.2339584, 1.2406066, -2.4173416, 0.0670238, -0.6658832, -1.8936084, 1.8712392, 1.6500735, -1.4947189, -2.0133758, -0.2487310, -1.4736210, 1.8683703, -1.2057520, 0.8722299, 0.3822608, -1.0009790, -0.4047141, 2.8308589, 0.4101696, -2.6062784, -2.5249203, 2.2124099, 2.7481077, 1.9686261, -2.5630033, -0.0470647, 0.6906985, -2.9218162, 2.2342638, -2.2415202, -1.2457207, 2.3692787, -1.9072749, -1.6720168, 2.9398599, 1.5313638, -1.7368440, -0.8653670, -2.8667395, -2.2368377, 1.5672557, -0.9745371, 2.4318524, 2.0896633, -2.2249317, 2.8470985, 1.5094681, 2.5866131, 2.0977633, 0.4158528, 0.6868469, -1.0133203, 1.2438762, 0.2674481, 2.5554143, 2.5111435, -2.4583223, -0.5512850, -1.2671767, -0.2448031, 2.0126427, 1.1948219, -1.8506911, -2.5532227, 2.5534149, 0.6201944, 1.5681238, -1.7962979, -1.9182889, -0.3100005, -0.2471829, 0.1456644, 0.8864958, 2.3187618, 1.4595516, -0.5172049, -1.1797177, -1.7064196, -2.1625613, 0.8653887, 0.9380741, 1.9001369, 0.3492953, -2.1708560, 0.4670710, -0.5072337, 1.5550823, 2.1141210, 1.9352925, -2.4414765, 1.8098044, -0.1984258, 0.2049534, -1.7574825, 0.5067826, 0.2732046, 1.9687988, -0.3706300, -1.1022542, 2.7107163, -0.8558547, 1.5408489, 1.8202093, 1.8991653, -0.8106989, 1.5243197, -2.6285289, 2.0085198, -2.7185629, -1.0124019, 2.9605110, -1.0569486, 1.5337522, 0.3602249, 0.0825543, -2.1801928, 0.1141204, -2.0723797, -0.8502576, -1.6922622, -0.1702874, 0.3199613, 2.6662362, -2.9178703, 1.2091079, -1.7031453, 0.6169439, -1.5381192, 2.3492964, 2.6655148, 0.2140390, -0.9962552, -1.6617311, 2.2131925, -1.7759480, 0.2228317, 1.4959877, -0.1305676, -1.3088267, -2.6882012, 2.6726292, -1.5957320, 2.8072158, 0.4961235, 2.6082411, -2.2333234, -0.5287335, -1.0173511, -2.7934046, 0.9941222, -1.7887470, -0.1980046, -1.4132971, 1.5244776, -2.0244737, 0.4828311, -0.3332968, -1.1254342, 2.6925746, -0.3462526, -0.9776232, -0.3318066, 1.2652640, 1.1566908, -1.0438177, -2.5299683, -2.8737725, -0.3177188, -2.0871784, 0.2473391, 0.5677394, -1.0803010, 1.7532660, 1.3586642, -2.9293779, -2.7880706, -1.5691156, 0.5159640, 1.9442837, -1.5276202, 2.4389329, 1.3383737, -2.0545479, -0.6761466, 1.6883263, -1.5670188, 0.1998539, -0.7595033, 0.2879874, -1.3016703, 1.4068899, -0.3046499, 2.9685089, 0.4771452, -2.2538908, 0.8325124, 1.0435475, -0.6534860, 2.3515131, -1.9515963, -2.3089604, 1.8942842, 1.3812240, 0.2831622, 0.6621886, 1.2152997, 1.6755728, 2.7885925, 0.6437487, 0.1334530, 0.1164920, 1.5479849, 1.7786499, -2.9434660, -0.2426165, 2.5371168, 1.1276626, -1.8337541, 0.4142883, 0.2236996, 0.3811593, -2.2475616, 2.0821669, 1.9103124, -0.8653258, 1.4176510, -2.7793514, -0.3602809, -0.3720276, 0.5531943, -0.0842706, -2.2168013, -2.2510958, 1.9742632, 0.3888652, -1.4182786, -0.5055101, -1.7738772, 0.0647455, -2.1427792, 1.7257930, -2.2803527, -2.8522793, 2.1577665, 0.5839522, -0.0338891, -1.1311412, 2.3110290, -1.8185918, 0.7141840, -1.0646775, 1.8510561, -2.0505600, 0.0669598, 2.1521601, -2.4754850, -0.3828349, -1.8745252, 2.4408168, -2.8953428, 2.8853897, 1.1984867, 0.2642965, 1.1327758, -1.8306042, -1.0020624, 0.5299732, -1.5225439, 1.3815068, 0.4910743, 0.5185269, 2.0280579, -0.9811543, 1.9192356, -1.4636742, 2.9862406, 2.6791544, -0.7066888, 0.6106749, 1.4788169, 2.9967702, -1.3928860, -2.9203479, -1.3170602, -0.9299529, -0.7652835, 2.4786277, 1.2923887, -0.3340939, 0.6905432, -1.6395410, 1.1220899, 2.0695880, -0.3684810, -1.7853020, -2.8752222, -1.7597800, -2.7739173, -2.4716397, 2.4808518, -1.0802492, 2.6777066, -0.0816514, -1.1222697, 0.0711571, -0.0923167, -1.1108268, 1.2292386, 1.9916046, 1.2506787, -2.0034849, 0.4190740, 1.9811586, -2.9710360, 1.9105262, -2.3341597, 1.6639581, 2.8882213, 1.4471022, 1.2311703, -0.7445011, -2.0809042, -0.2180699, 0.8479292, -2.2911788, -0.1192878, 0.1204366, -1.9824434, -0.5443266, -1.7350627, -0.5310373, -2.1971262, 2.3610731, -1.5689469, 2.9795764, 0.9431471, -0.9781985, 2.2033260, 0.8735649, 2.3835714, 2.3415948, -0.8808307, -0.7057753, -0.9402073, 2.7965031, 2.8844060, -0.8401587, 1.3594178, 2.6540376, -1.9664905, 2.3889390, 1.3579128, -2.7227150, 1.6401132, 2.5165632, -0.9105365, 2.4721122, -1.1953450, 1.4231590, 0.3414116, 2.3000166, 2.1616719, 0.0025036, -2.8472292, -0.0743712, -1.8083889, -0.0068304, 1.4075656, 0.2823809, 2.3592689, -2.8075985, 0.8125600, -2.6427540, -2.4029534, -2.7832333, 2.9337061, 2.1503571, 0.2346175, 1.7595205, -2.4372863, -1.3804633, 1.2830502, 0.4793136, -1.3443367, 2.0424424, -0.0747316, -0.8706969, 0.2177267, 0.1136518, -1.0425937, -0.6596061, 2.7151037, -2.8542585, -0.7734686, 0.6824353, 1.0161111, 0.2746939, -1.2428468, 2.2598531, -1.2049485, 0.2175512, -2.4815444, -2.9417080, 2.8853870, 2.2636913, 2.2464362, -1.4306303, 2.6256221, 2.6206791, -1.1610948, -1.1703297, -2.9220676, 0.9526531, 2.3178087, -0.3903316, 2.1875056, -0.4301841, 1.1615198, -0.0038952, -1.5525895, 2.2817627, 2.7717375, -1.2160243, -0.0369598, 2.2046336, -2.1172752, 1.4305392, -2.9958612, 2.8843682, 1.0157875, -0.4525454, -1.1391363, -2.3658554, 1.7235305, 1.7131144, -2.9470302, 2.3286755, -0.7310478, -0.2175845, -0.5326366, -2.2340692, 1.1707722, 2.6033538, 2.6102216, 1.6295904, 0.3227767, 0.6733060, -0.0958410, 1.8534636, -1.6265420, -2.4119545, -2.1419230, 0.4339400, 2.9957601, 2.9574385, 0.6903105, -1.6082384, 1.1111469, 0.3869265, -2.1358842, 1.1851412, -2.4095148, -0.2456741, -2.9718662, 1.8014557, -1.4850717, 0.5121619, -0.8237835, -1.9493982, -0.4027002, 1.5898046, -0.6019064, -0.6865683, -1.3297408, -2.2841372, -0.9130129, -2.7425367, 1.9831361, -0.7270325, 0.0689664, -0.7754405, -2.3691769, -2.7427054, 2.3703015, -1.5585993, -1.5963479, 1.7501044, 2.3117388, -1.9086453, -2.3496304, -2.6812473, -2.7282186, -0.7857225, 0.4626504, -0.5920170, 1.4118287, -0.9067660, -2.7037969, 2.1528972, -2.7614172, 2.2135483, -2.8035996, 0.3584441, 0.1450736, -2.7715720, -0.3858994, -0.4046132, 2.4899711, -0.2039436, -0.1608280, -0.8519998, -2.8316055, -2.9159462, -0.3898225, -2.1538384, -1.6193002, -0.3725714, 2.6007230, -2.6677293, -0.3919114, -2.0265986, 0.7924420, 0.4016495, 2.3478331, -2.0962630, -0.8043476, 0.5695782, 2.9488293, 0.8249305, -1.2033894, -1.7122684, 2.4030487, -0.4656143, 0.1244416, 0.9944613, 0.6246107, -0.7784354, 2.5379289, -2.8974280, 0.0092865, 2.5366995, 1.8490610, -1.1738958, 2.7010514, 2.3720957, -2.8600192, -0.5120816, 0.4523638, 2.2248258, 2.6955626, -1.5104240, 0.4065943, -2.2618674, 1.1084334, 2.4029223, -0.4931995, 1.5203954, -0.2087817, -0.6641746, 2.6070881, -1.6925528, 0.3658673, -2.1631240, -2.1395142, 2.5180269, -1.8220605, 2.7296194, 1.6401129, -0.7053914, 0.6239152, 2.1744587, -2.6812658, 2.5787870, -0.1044783, 0.0897259, -2.7724836, -1.1877838, 1.0849980, 0.8763878, 1.7064406, 0.7915039, -1.5818355, -2.9407369, 2.0299960, -0.3196668, 2.3360228, -1.8956208, 2.0285027, -2.9055316, -1.8367038, -2.0101763, -2.1463051, 2.5080507, -0.4291403, 1.1951042, -0.7449050, 0.7077184, 1.0252296, -2.9169975, 1.6509952, -0.4829813, 2.7792818, 0.2479234, -2.4434816, 2.0499442, 0.0000149, 1.9159751, 2.5375098, 2.4621610, -0.8993375, 1.5970055, 0.8552119, 2.8793330, -2.1884453, -0.9076832, 1.7603060, 0.0488743, 2.7457980, 0.2150499, -1.3281986, 2.7368659, 1.6537978, -1.1121448, 2.0894953, 0.7534505, 0.2311128, 0.0697528, 2.8148851, -2.6193658, 0.6391138, 0.4143829, 0.1297927, -0.0659273, -1.4423078, -1.6648113, -0.0678345, -2.8022935, -1.8484089, 2.3960694, -0.3153642, 0.1136888, 2.6517462, -1.8444899, -0.7150561, -1.7343226, -1.8667321, 1.7315830, -2.0238566, -1.9769380, 0.5827283, 0.2783295, -2.1203601, 0.0782977, -0.6956679, -1.8376185, -2.5758577, 1.8667640, -0.9971535, 2.8131011, 2.9783418, -2.8751351, 2.0519444, 2.7500878, -1.5695240, 2.6817346, -2.0109634, 1.8290616, -1.6551013, -0.4779843, -0.0981002, -1.7056951, 2.4693347, -0.2931356, -0.9781127, 1.5631455, 1.8173530, 2.5747959, 2.3221010, -1.1928952, -2.8494765, 2.2720845, 0.7045294, 1.9331593, 0.9558378, 0.0415443, -0.7035737, 2.1454370, 1.5155774, 1.1820183, -1.1966597, -1.8842746, -1.1444680, 2.1482492, -1.7158941, -2.0364947, -2.9809163, 1.4161161, -1.4261547, 0.2801366, 0.2494508, -0.7355653, 1.2960990, 1.3503174, -2.4847039, -0.2588250, 0.9138741, 0.1682822, 1.0939725, -2.7372736, -0.8332990, 2.9055581, 0.1824591, -2.2837603, 2.1075854, 2.4591047, -2.1174846, 0.0140805, 1.5625309, 1.5189219, 1.2311848, -2.5107199, 0.4880808, 2.3191603, 1.9969393, -1.0349719, 2.9790860, 1.5231985, -2.0541559, 0.1257887, 1.6568434, -0.5747511, -2.6248384, 1.0326363, -0.7130838, 1.2719305, -2.0676256, 2.9866839, -0.6313003, 2.0202651, 0.3492021, 0.5263524, 0.5390430, -0.0940016, 1.5884298, 2.7364612, 1.6585858, -0.5927766, 0.8975355, 2.7092084, -0.6236759, 2.3285204, -1.1568772, -2.7698510, -1.5730351, -0.5509250, -1.5975664, -2.0302069, 1.1990098, 1.5155930, 1.6948288, 1.7610739, -2.7681563, 1.3253927, -2.4002901, 2.5212613, 0.8958430, -1.3149503, 0.8691733, -1.6360879, -1.9906013, 1.9209638, 2.0330408, -2.9847171, 2.4661194, 2.4412083, -2.8157749, -0.8237896, 1.6956267, 0.7415755, -2.3018833, -1.4269063, -1.0934620, -1.5786555, 2.3720534, -2.7393565, 0.5616599, -0.4828762, 0.2450424, 1.0682854, -2.7007128, 0.9574407, 2.3503262, 0.0500976, -1.8461306, 1.1200064, -1.0389711, -2.9388277, 0.5527264, -0.1642845, -1.3592605, -1.7351357, 2.2903713, -1.6318264, 1.7351670, -1.6951667, -1.0437263, -1.4323671, -2.4633894, -0.3326340, -1.3352984, -2.3287763, 2.6773888, -1.5414750, -0.4974105, -0.5260775, -0.1020058, 2.4654978, 1.5072612, -1.8145679, 0.7771501, -0.5148989, 2.6461342, 1.5855155, -0.7397477, 0.8389943, -0.9526401, -2.4906874, -0.2407649, 1.7919140, -2.4687487, 0.7206562, -1.1202191, -1.3528318, 1.7466294, -0.7280075, -0.0490011, -1.7971141, 0.0959833, 1.2553179, -2.8983254, 0.5772709, -1.8705179, 0.2253020, -1.5726284, 1.8704064, -1.4423504, -2.3729368, -1.1257585, 1.5989019, 2.9820202, -1.3212801, 1.5956682, 1.7299917, 1.8686605, -1.2913184, 0.5478053, -0.1664510, -0.7342943, -0.6402617, 1.8271064, -0.5671919, -2.0708659, 0.6570476, 2.1867386, 0.0241932, 0.4880007, -2.3293203, -1.1911982, 2.3927353, -2.1081908, -2.6062009, 2.5403035, -2.9006758, 2.4938934, -2.3259367, -1.4179663, -2.2201298, -1.2700978, -0.4720458, 1.8157385, 0.9780604, -1.6583172, 2.3659216, 2.5712648, 0.9184561, 0.0788216, -0.0408175, -1.5650978, 0.5363412, 1.8437786, -2.7667762, 0.5204136, 0.8529482, 0.0439042, 2.9252867, 2.2470342, 1.7452539, 0.8222188, 2.6050044, -2.4780261, 1.4124408, 1.4833955, 2.0135334, 2.8002818, -2.3786086, 0.9269775, -0.6407230, 2.5437605, -0.6451810, -1.4873298, -2.5984053, 2.1976952, -2.2965321, 1.6555807, 2.4311753, -0.8177269, -0.9243594, 2.8418836, -0.0988785, -1.3474955, -1.8993681, -0.2163328, 1.7717038, 2.8693233, 0.6223830, 0.3827387, -1.3754498, -1.0061520, -0.3524990, 1.3790492, -2.4548934, -0.8689708, -2.0452031, -1.5082795, 0.4212828, -2.0875795, 1.7419588, -0.7260314, -0.5371284, 2.1923640, -2.7666701, -2.6844846, 2.2813021, -1.3942406, -1.3867380, -2.7828333, -2.1158219, 1.9725495, 0.4847222, 2.4132298, -0.8795818, 1.1759323, 1.2586685, 2.2196521, -2.5586607, 2.4594953, -2.0305114, 2.8766704, 1.7323006, 0.7693855, 2.6046159, -2.2849192, 2.3749248, -2.5865987, 2.6056384, 1.5587254, -0.9249990, -2.7167961, -2.1461192, 0.6672778, -2.9194273, -1.5111461, -1.2356426, -1.5997979, -0.1490678, 0.6719964, 1.0651910, 2.8591804, 0.9369508, -0.9846423, 0.0437022, -0.8343176, -2.5210329, -0.4052211, 2.8969494, -0.8066030, 0.3939007, 2.2999768, -1.4112426, -1.5422073, 1.7404740, 1.6800065, 0.5374487, -1.7692288, 0.9008447, -0.8976867, -1.0605374, -0.8312649, 0.7492257, 2.0845628, 2.7985147, -2.1869561, -2.0803345, -2.1064283, 2.1598971, -0.6036671, -0.7033672, -1.0377670, 0.5670020, 0.8397677, 1.2562394, 1.9809762, -2.6740966, 1.5598853, 2.3746351, -2.6380644, 0.6484097, 0.3152243, 1.1513564, -0.9003889, 0.7519242, 1.6231223, -1.1339935, -2.0922143, -1.9091807, -2.7191499, -0.6449160, 1.1810213, -0.0584696, 2.6441348, 0.4401933, 0.6717545, 2.1241526, 2.5018782, 1.4501555, 0.2445915, -0.9787351, -0.6706115, 1.9913328, 2.1131990, -2.5983321, 1.9173641, -2.8320931, 0.7788981, -2.8602817, 1.5985833, -2.3162411, 0.9011583, 0.7996340, -1.4896151, 1.8601751, -2.9016261, 2.3007984, 1.9402835, -0.1281197, 1.4557902, 1.0449109, -1.0010384, -2.2043371, -1.9212375, -2.5192120, 2.7433096, -2.6189941, -2.5451047, -0.1819037, -1.1774380, -0.3684874, -0.1398540, -1.4096586, 1.7783095, -2.0731444, 0.5067611, 2.6206657, 0.5321105, -1.1597214, -2.0239307, -0.3169768, 1.1385887, 0.6278899, -2.6174629, 0.9312676, -0.3168756, 0.5970354, -1.0124716, 2.5072666, -2.0121583, -1.7039640, -0.6121936, -1.1124305, -0.6244704, 1.4982441, 0.5025140, 0.8831703, 1.7339467, 2.7217198, 1.7840383, -1.4402152, 1.6497295, 2.7702613, -1.0464755, -0.1480127, 0.5340051, -0.4662509, 1.3178280, 0.4208277, -1.5860057, 1.0029543, -1.6074332, 1.0117810, 1.2094674, 1.1914707, -0.9364509, 2.1107302, 2.3745303, 0.5595874, 1.1545669, -1.0789893, -1.5690228, -1.9867564, -0.6642873, 0.8452624, 0.9937033, 0.1734226, -2.0883607, -0.9104947, -1.6543876, 0.5314960, 1.4218704, -0.4548378, 1.3654905, -0.7682956, -2.0426459, 2.0659442, -1.4139894, 2.2101927, -0.4944643, -1.5608702, 2.2961658, -2.9575702, 0.5760243, 2.8364763, 2.3312013, 1.0579933, -2.3591658, 1.3387576, 0.3634454, -2.6687960, -0.5265401, 1.8445088, 2.4203792, -2.5806122, -1.0897797, 2.3111960, 0.9922565, 0.6375720, 2.8382158, -0.8154290, -1.0552812, 0.7277475, 0.9541958, 1.7363045, -2.0448585, -0.9152923, -1.7443739, 1.8015563, -0.3278642, -1.8867711, 1.9503284, 2.1532829, -0.7854651, 2.6752043, -1.0875309, -1.6556629, 2.8239888, 2.1344657, 0.8737221, 0.8388017, 2.4738452, -0.3582608, 0.5595618, 1.9715996, -0.0827810, -2.2100553, 0.6428994, 0.0714283, -0.5859359, 0.2070983, -0.0769194, -2.0073572, -2.4236956, -0.2475665, 1.5650586, 1.4787881, 0.8371356, -1.9056666, 1.7814827, -1.0550810, -2.4583902, -1.2674971, 0.6484995, -1.5987224, -1.0942791, 0.0347767, -1.2916928, 2.1040917, 1.5689450, -0.6157620, 2.8095943, 1.4431533, 2.5407794, -2.6660289, 2.0481999, -1.5758322, 0.9040177, -2.2938788, 0.0133825, -1.3597069, 1.3466394, -1.5319545, 2.7369299, 2.1924768, 0.5312385, -0.2781351, -0.3695590, 2.2769142, 2.7050995, 1.6819414, 0.8124177, 1.3976342, -0.9156871, -2.9389622, 1.0624109, -0.2668143, -0.1023114, 0.8274295, -1.3635918, 1.5715082, 1.5664033, -2.7805803, 1.7876932, -1.9416154, -1.6747901, 0.7921690, -2.3356901, -0.8419595, -2.7765363, -2.9850564, 1.5768317, 1.4350734, -0.9029670, 2.5093045, -2.0753570, 0.6343162, 0.6066664, -1.9104795, 2.2972883, 1.7871607, -0.4561123, 2.0882792, 0.6132840, 2.9327215, 1.5553455, -1.0505546, 2.8593854, -2.3230401, 1.0280402, 2.8265192, 2.7380527, -0.8639773, -2.6318872, 0.5310477, -2.6661619, -0.7556020, -0.9733746, 1.3792919, 0.6187133, 0.8068820, -1.7675950, -0.8083932, 2.9139210, -2.5070434, 1.6824209, -2.5288309, -1.6929706, 2.0681442, -0.2806894, -2.7900149, -0.3207714, -0.4618045, -0.5450293, 1.8971913, -1.7962719, 1.3182918, 1.2531096, -2.2659037, 0.4671628, 0.9229102, 1.5158068, -0.4233742, -1.5171685, -0.5885423, -0.0340415, 2.9297989, -2.3322490, -0.8434190, -0.5988848, 2.1848315, -1.8439187, 2.1147281, -2.5798434, -2.2286576, 0.7220271, -2.8975673, -2.2005381, 0.5222942, -0.3677996, 1.5886045, -0.5335281, -0.3026308, -0.8894725, -0.3267679, 2.0940960, 1.9932741, 2.9216625, 1.0759281, 0.0209866, 0.1454837, -1.0511640, -0.5683806, -2.2382295, -1.3118743, -1.7179858, -0.7084533, -0.2892322, 0.0492360, -0.2533827, 0.1040820, 0.2567953, -1.2523362, -1.6016147, -2.9515425, -0.7054476, 1.8117171, -2.9366680, 0.7544765, -0.1191087, 2.1113413, 2.6540952, 2.3678368, -1.7594267, -0.0281247, 2.2390566, 2.3867173, -2.4680441, -0.2561858, -2.4383062, 0.7716993, -0.3973376, -2.0866204, 0.4463396, -0.6041492, 0.4245564, 2.5172230, 2.6268425, -2.1752439, 1.7152455, 0.3961999, -2.4742472, 0.9647532, -2.5456254, -0.2231310, -0.9530808, 0.1622072, 0.9398284, -1.0875351, 0.3070245, 0.3774869, -2.8623201, 2.0360449, 1.8908233, -2.4188701, 2.4863789, 0.9747363, -2.6644412, -1.1856047, 2.4349155, 1.4438559, -2.9278715, -2.3027470, 1.9405459, -0.2833653, 0.3887457, -0.1421806, 1.6119555, -0.9795003, 0.6556764, -2.5063434, 2.7038403, -0.1021164, 1.1514915, -1.6962669, 1.8985263, 2.7816922, -1.0240801, -1.3916377, 0.1351129, -0.6765417, -1.1946720, 1.5679435, 1.9202122, 1.1109269, -1.9388213, 1.7801632, -0.2940811, -0.4354091, 0.9575495, -0.6545514, -2.5501337, 1.5384968, -0.0443361, 2.1507623, 0.3918269, 2.1392035, -0.4339557, -2.0333465, 1.8751724, 0.7987049, -0.8531825, -0.4784860, -0.6277742, -0.2648143, 1.7975673, -2.4503609, 1.3578642, -1.6598590, -1.7294517, 2.8556123, 2.4073585, 2.7497366, 0.8531307, 0.9370011, 0.3161322, -2.7874382, 1.3258935, 0.3860629, -1.4630127, -1.1951268, -2.3533152, 1.8416516, -1.3590486, 2.3147601, -0.0264726, -1.9755962, 1.3495156, 1.1212933, -0.0263620, -1.6314486, 0.4719112, 0.6984047, -2.3275829, -2.8919267, -0.7635236, -0.9341350, -1.9954382, 1.2278332, -2.5223434, -1.5444316, 2.2471759, 0.8927175, -1.2601156, -2.7249806, 1.4087667, -1.7773878, -0.4759638, -0.9579910, -0.7109819, 2.3555727, -2.8940594, 1.3389484, 2.1832813, 1.5158027, 1.2436744, 0.4665205, -0.6326685, -0.4258846, 0.7626476, -1.8286210, 0.5610973, -0.7811548, 2.3178142, 2.6889441, 1.7163479, -2.3788704, 2.9115103, -1.2953107, 1.5700387, -0.2582557, -1.9783932, 0.3479013, 2.6153557, 2.0354347, 0.9645193, -0.3645705, 1.0901428, 0.8825376, 0.2363209, 1.6869969, 0.7481373, -0.6433627, 0.6962408, -2.0067565, -2.6071389, -1.7011510, -1.3964278, 2.6058783, -1.6300902, -1.1089887, -2.7693138, -0.0228391, -2.5716231, -0.9057979, -2.7851950, 2.6556163, -2.0351794, 1.0822693, 0.4305640, -0.9119288, 2.1732969, -0.2108484, 0.6911821, 2.6570519, 2.1352629, -0.9275853, -1.6642185, 2.7535613, -2.3064658, -2.8174513, 0.3383563, 2.4341015, -0.2581573, 2.2287009, -2.5026158, -1.2168167, -2.8368007, -2.5724502, -2.4103078, 1.1842593, 0.1648137, 1.1284911, 2.8200416, -1.7411088, -1.1121489, -2.0895377, 2.3540753, -1.9114320, 0.4427727, 2.1182141, 0.0610017, 2.6869325, -0.9349935, 1.2273653, 1.6178831, -2.2668077, 1.0180328, 2.9471954, 0.7873251, -0.9214316, 1.0760165, -1.0217538, -0.6935015, 2.0555052, 0.8202207, 2.5370686, -1.1903733, 0.7282211, -2.6359046, 1.7224118, -1.4308375, 0.5021813, -1.5938267, -2.5503764, -0.5722040, 1.7947884, -1.4836415, -2.9222332, 2.2437798, -0.7369683, -0.1061404, -0.5956211, 1.8108897, -2.3189248, -2.9669738, -1.8143315, 0.3504712, 0.1015704, -1.0587351, 0.1255807, 1.7926296, 2.1299803, 1.4655581, 2.2330186, 2.2883719, 1.4818756, -0.3634864, -0.0872399, -0.4061504, -1.9599298, -1.4613517, 1.1288030, -1.0974817, 2.1507981, -2.6587974, 2.1478687, 2.2431260, -2.5577244, -2.1415483, -1.3249047, -0.7808485, 1.5992910, -0.5781948, -2.3537064, 1.9997751, -0.0563151, 0.0675561, -2.2381240, 1.6465217, -1.1229448, 2.3856507, -0.8545700, 0.6569760, 0.6402804, 0.7723737, -2.1745804, -2.6946882, -1.6373203, -2.2498785, 2.3622937, -0.6200435, -0.4237836, -1.5541667, 2.3277666, 0.2663014, -2.5328250, 1.0951499, 2.8334155, -2.4399769, -1.2616428, 2.7603339, -0.4678929, 1.7191764, 2.9564476, 1.5576801, 0.0345115, -2.6194780, -0.0247523, -1.8875676, 2.0541651, -2.6818356, 2.8257374, -2.7909271, 0.8470850, -0.9414999, -2.6336532, -1.9866870, -2.0381695, -1.3864981, -0.2703132, -2.2183736, 2.7604007, 2.9002182, -1.0384397, -0.8615894, -1.6022648, 2.9651349, -2.0367814, -2.3047264, -0.0449928, 0.6152981, 2.6513565, 2.7324473, -2.3914379, -0.0174146, 2.6694070, -2.0441010, -2.1250370, -2.1604680, 1.5686897, -1.5892230, -1.7291031, -2.2290314, 0.7162180, -2.6345731, 2.1671987, 0.4951155, -1.8523150, 2.5306053, 0.9836286, 0.8152677, -2.2104383, 1.0611336, 2.1947311, -2.4922968, -1.3680954, -1.4280416, 0.2997870, -1.7375998, -2.2041637, -0.3971372, -2.1327234, 2.2190545, -2.3376279, 2.2431574, -0.5781253, 1.8307615, -0.3894057, 2.0316595, 1.7770613, -2.2113781, -0.8743625, -1.0671462, 0.8235078, -0.7273056, -2.9561605, 0.9602164, 0.7893213, 0.8252352, -1.4239553, -0.4330352, 2.9731040, -1.8903038, 0.0187190, -1.8321509, -1.7845871, 2.2735606, 2.0715570, -0.7711800, 1.3480032, 0.9825389, -0.3343296, -2.8148937, 2.2097089, 0.0685234, 2.9240478, 1.7932637, 1.9800566, -2.1720415, -2.0083751, -2.2915463, 0.5315251, 0.3991659, -1.9014110, 0.2038770, 1.2667053, 1.0770633, -0.9076861, -2.3091168, -0.8060541, -0.1287503, 2.9659467, 1.7362288, 1.7907845, 0.2964916, 1.1402125, -1.3663742, 2.5099394, 1.6033162, -0.7550353, -1.9445734, 1.3216664, 2.8881317, -2.0391145, 0.7337443, 0.4542729, 2.6157209, 1.5095767, -1.9394514, 0.3981010, -0.7548715, -1.7788062, -2.4762798, -1.7585121, 0.2513674, 1.3138048, -0.4239607, 2.7377924, 2.1521100, -0.4594306, -0.6634807, -2.5911153, -2.2653204, 2.5028556, -2.5304333, 1.8288843, -1.5675195, -2.8833131, -0.4180928, -1.3628700, 2.1779490, 2.4567891, 2.4244278, -0.5622605, 2.9662835, -2.0836879, -1.0860557, 1.9893431, 1.2940240, 1.0475765, -0.1382839, 2.0138845, -0.9093208, -1.0065755, -0.2485959, 2.2458792, 1.7969524, -1.5207555, -1.3300628, -2.1087579, 1.4106679, -1.4582444, -0.8285658, 0.3042878, -2.6589236, 0.9564894, 0.3339710, -1.4383295, -0.9560151, -1.5086579, -2.3349462, 2.4294745, 0.1937332, 0.6443203, -2.9290670, 0.1954825, -0.9796684, 2.7305542, 2.2271710, -2.2445970, 2.7173397, 0.6041717, -1.4100180, 0.9219241, -2.7903708, 1.6914851, -1.7409681, -1.8614774, -1.0895926, 2.3011757, -1.1508175, -1.4176801, 1.3726045, 1.2292122, -1.8576230, -1.4233208, -2.0664593, 1.8919352, 2.1343955, -1.5120053, -2.1012035, -1.6433305, 1.1505144, 0.8863140, -2.2484079, -2.7610188, 0.8311473, -2.9807737, 1.3819376, 1.2372104, -1.0729090, -1.8779353, 2.7689559, -0.4813131, 2.8078546, 0.0336725, 1.5360088, 0.4999941, 0.4383989, 0.5482611, 0.6852272, 2.8652333, -0.6805215, -1.4557755, -1.5856394, -2.5073283, 1.5981613, 2.8791269, -2.9611676, -1.7452746, 2.3976670, 0.5217198, -1.0915379, 1.2854252, 2.7158146, -1.5486111, 1.0405933, 1.2887423, 2.6010468, 0.4638997, 0.9150854, 1.0867427, -0.8971788, 0.2512148, 0.3069637, 0.2689059, 0.1790002, 2.1662842, 2.9280104, 2.8107625, -0.6843840, 2.3262566, -1.8779674, -0.4555090, -0.7055956, -0.0852931, 1.5855352, -0.7040596, -0.3483318, -0.8484567, 0.2853106, 0.2066325, 2.5175130, 1.7347753, 1.8647922, -0.7897539, -2.1164916, 1.4330947, -2.3734319, -0.3457963, -0.4505273, 0.6692436, 1.6799523, -0.9154607, -1.2613139, -1.6077096, -2.6902363, 2.5084108, 0.1793430, -1.9340245, 1.5662247, 2.0923664, 2.0360888, 2.9212474, 2.0045283, 0.3658087, -0.7004799, -2.6553424, -1.8619484, -2.1353143, -1.9911259, -0.2414117, 2.9453189, -2.6643556, 2.6536626, 0.9123664, 0.1431236, 1.1932030, -2.3256796, -1.5133548, -0.0541543, 1.4003426, -0.1451357, -0.1472083, 0.3524763, 0.8554287, -0.7955038, 1.7017694, 2.5848436, 2.8468825, 1.8623698, 1.7325561, 2.2389634, -0.6878645, 1.8270873, 0.0738046, -2.4091611, -2.0965360, -2.7244852, 0.0000447, 0.6623941, 1.7243674, 2.2701985, 1.2824159, 1.3173242, 0.3396739, 2.3699363, 2.4376645, 0.9773146, 2.0470504, 2.6182562, 1.5048674, -2.8072625, -2.5058078, -0.7302034, 0.2135305, 1.2113683, 1.6880778, 0.1942946, 2.2753237, -2.3644032, 2.6829166, 2.5445571, 0.1412452, 0.2272834, -2.7087310, 0.8463212, -1.2377812, -2.2975514, 1.3452304, -0.3108132, -0.4526783, 1.4080700, -0.3668269, 0.3098688, 2.6996596, 0.6147868, -1.7258265, 0.2077745, -0.3037452, -2.7858178, -1.1098688, -2.2011803, 2.9973158, -2.7640046, 2.9987602, -0.0683403, 2.0897097, 1.2818047, -1.1589155, -0.7990811, 1.7823346, -1.9223970, 2.5985602, 0.4455628, -0.8434308, 1.3811717, -1.9941865, 0.8644776, 1.8467580, -1.8339982, 0.3411223, 2.8489680, -2.9330269, -2.7871312, -0.5986596, 0.3791222, -0.3781309, 2.0876544, -1.5070658, 2.7066606, -2.5607881, 0.2100686, -1.3680852, 2.7733853, -2.3266224, -0.5510000, 1.5456266, -1.5156962, 0.3338931, -0.5958959, 2.0496420, 1.8383114, 1.8877420, 2.9040294, 1.9201950, 0.4490231, 2.0416814, 2.6389264, 2.7664695, -1.5752078, 1.4323611, -0.1102555, -2.1393119, -1.7902889, 2.1468586, -2.0123684, 1.7307831, 2.8976087, 1.3063662, -0.6726304, 2.4200498, -2.1456511, -1.6996109, 1.1025184, 2.8357695, 0.4834362, 1.0233508, -1.2473967, -1.0777573, 0.2804416, -1.9942486, -0.9913350, 2.1220607, -2.7756803, -2.0250503, 2.9548878, 1.3760192, 1.8547075, -1.4688001, -0.4482630, -2.7706386, 1.7466239, 1.1632696, -2.9848459, 1.3427539, -0.9662957, -0.8516734, -1.6765704, 2.0344362, 2.6362304, 1.1106716, 0.5802483, -2.6203796, -0.8070918, 0.1719766, -2.1458403, 0.1324252, -1.1933531, -2.5029833, 1.8284851, -1.9059811, 2.0699075, 2.5829430, 2.2749770, -2.0862537, -1.3261655, -1.7640727, 1.4152452, 0.0058173, 2.5379568, -0.4815041, 0.1768406, 1.6237120, 0.9806167, -0.5320896, -0.9376097, 2.7628802, 2.2872849, 2.4929525, 2.4741022, -0.5990682, 0.0450778, 1.5358188, -0.1537173, -0.9141683, 2.9685662, -2.0094547, 1.3916661, -0.8909597, -0.5822857, 1.5623925, 0.4062776, 0.4762293, -2.3096791, -2.9084707, 2.9027549, -2.0982564, -1.5135441, -0.3606733, 0.5027039, -0.3669662, -1.3711208, 0.5910628, -2.0102363, 0.4305492, 0.4196680, -2.5605661, -0.6154318, 2.8832469, 2.3691537, -2.3643376, -0.3028799, -0.7818446, 0.8667011, -0.1686067, -0.1257021, -1.0119683, -1.6095102, 1.7046300, 2.8770683, 2.2123770, 2.3059197, 2.7685406, -1.0789232, 2.3722002, -1.0684453, -0.8944371, 2.5535144, -1.6640974, -2.8219046, -1.0363543, -1.3607160, 2.0605889, 0.6527418, 0.6051551, -2.9434803, 1.1019667, 0.4307406, 1.4712792, 0.6900596, -2.3476424, -2.9757350, 0.8819655, -2.6815447, 0.9897053, 0.7106965, 0.4403465, 0.1980361, -1.9849771, 0.3204066, 1.2785296, -2.5618454, 0.2802101, -0.5546306, -2.3712417, -1.5285317, -1.1931052, 1.2129608, -1.2108811, -0.7529158, -1.1893094, 1.0457340, -2.9226409, -0.5899036, 1.7368112, -1.5016926, 2.6136037, -0.6679030, -1.9096958, 2.3056247, -2.8711132, 2.6578285, 1.6401000, -1.1624869, -0.3543876, 2.5957145, -1.0203609, 0.5869389, 0.1650516, -0.1878482, -2.4274901, -2.2540330, -2.5072510, -0.7987803, -2.0385402, 2.7926004, 1.6968126, -0.2058793, -1.0053841, 2.5155506, -2.7519839, 2.9730731, -0.4000398, 1.0434298, -1.1825903, -2.4276836, 0.1174220, -2.4691665, 1.7050402, 2.8695352, -0.1659990, -2.3702949, 0.5045314, 1.8153869, 0.7873690, -1.6119563, 1.7905436, -2.6474080, 2.9410395, -0.5849664, -1.6644115, 2.7149717, 1.9180602, 1.7881126, -2.4780497, 2.6105076, 1.9791806, 2.4098058, 0.1830881, 1.1075844, -1.7857334, -0.4366864, 1.9290081, -1.3355471, -0.4904798, 0.5805684, 1.4856772, -2.1306416, -2.6408679, 2.8690158, -1.7533735, -1.4071873, 0.5470582, 2.5191319, 0.4256519, -0.7979667, -0.3917049, -1.9471685, -1.9517761, 2.2017539, -1.1880746, -0.8841534, 0.1431945, 0.6977159, -1.8850628, -2.1396397, 1.2758792, -1.8603935, -0.9745877, 2.0431252, 1.3208626, -0.8998845, -0.2123021, 1.5501973, 0.8857457, 2.4895893, 0.7914235, -0.7901847, 0.0605593, 0.7467626, -2.2929315, -0.6514921, -2.4961831, 0.0112493, -2.5189143, 0.6277224, 1.6320823, 1.0912124, 0.1337701, -0.3416370, -2.1218108, -0.2508318, -0.4385385, -1.4148972, -1.7275931, -2.5016407, -0.1131272, 2.1372900, 0.1018040, -0.6732767, 0.8264508, -1.5983401, 2.9003362, 0.4406721, -0.0059236, -0.9604966, -2.9087285, 0.1140540, 2.5991266, 1.8141557, -1.6184122, 0.2326356, 2.2603501, 1.3502872, -0.6385021, -2.1896546, -0.5488877, 0.2147515, -0.0173332, -0.7411615, -1.0922811, -0.0587453, 1.9635825, -1.0675971, 1.3515601, 0.1408579, -0.5267947, 1.1002925, -0.1265364, 2.8050276, 2.9715413, -1.9568830, 2.1953545, 2.6718741, -2.9182236, -1.5845823, 2.5446625, -1.7670631, 2.8906762, 0.6926223, 1.3269907, 0.9783469, -0.9815578, 1.0657678, -0.1230469, -2.3729809, -2.3876580, -2.9317870, -1.7463910, -1.5783632, -2.4420435, 0.7577982, 2.4311502, 1.6186469, 0.9457338, -1.6472069, -0.3311809, 1.4051908, -1.1064961, -0.5239001, -0.1032929, -1.8264015, -0.8021071, 1.0914030, -1.1522563, 1.3115649, 0.5302698, 1.1322640, -0.3643352, -0.5340858, 0.8290348, 1.6289244, 2.1218302, 1.0537177, -0.5698514, 2.5552157, 2.1332736, -1.7106464, -0.3391859, -0.4495048, 0.7809156, -0.6967023, 1.7483999, 0.0950138, -0.9790270, -1.8014491, 2.8166342, -2.4252996, -1.5973610, 0.5575905, 1.0934681, 2.2009449, -0.7544189, 1.8591155, 0.6327589, -1.2847183, -2.2536194, 0.8036155, 2.3522052, -1.1391564, 2.2085496, 2.6443374, -2.6750020, 1.2319222, 1.0014629, 0.2805376, 1.6422078, 0.6529274, -1.8244049, -1.9700435, -0.8635928, 0.8759334, -2.7649350, 0.2751174, 2.8358570, -0.7788254, -0.9992282, -1.3776838, 1.7333980, 0.1739192, 2.1368746, 1.6544333, -2.7510212, -0.1632872, 1.2065347, -0.7753330, -0.1454972, 1.9064731, -0.6477096, -2.1048658, -0.3052030, -0.2576712, 2.7551546, 2.5938213, -1.8156483, -0.1414945, -1.3490267, 2.4238474, 0.4118564, 1.6454239, 2.6596310, -0.3066919, -1.0388598, 1.4949212, 2.1894232, -1.9008380, 2.0337884, -2.5724612, 0.2436428, -1.3386488, 2.2967611, -0.9358126, 1.6643984, -0.4868456, 1.2073076, -2.2636422, -0.2261495, 0.2654259, -1.9130571, -2.8453472, 0.5505948, 1.8191426, -1.8765364, 1.3755408, -1.4663266, -1.3268393, 2.3203500, 0.7058855, -2.9080440, -0.3794960, 0.6881935, -0.8580726, -2.5360564, -1.4008651, 1.0842597, 2.6716495, 0.8997241, -1.8569697, -1.8185107, 1.4640170, -2.7918926, -2.2176894, 1.7961929, 1.5042765, -1.2123884, -0.0598890, -0.3363615, 1.4358852, 0.0426488, -2.9014801, -2.1519741, -2.8511059, 0.7534012, -1.2723212, -2.5716095, -0.2931973, -2.6363919, -0.2295930, -0.5567242, -1.9254793, -0.1601815, 0.8330000, 2.8593257, -0.9515382, -0.5704676, -1.8057539, -0.7322481, -2.5383961, 2.7484140, 1.3963997, 2.9212113, -1.4306426, -2.7170233, 0.8440530, -1.0735038, -1.5694756, 1.6683532, -0.6531745, 2.9261031, -0.1741325, 2.6034237, 0.1939444, -1.8298936, 2.9975905, 0.4288863, 1.3076282, -2.0187927, -1.2393390, -2.4008633, -0.9114399, 2.7945251, -1.7679769, -0.0396249, 1.5348192, 0.3480056, -2.0980811, -0.1098128, -2.9094894, 2.3452192, 2.1023222, -2.8848616, 1.0966303, 1.3555133, -1.5083335, 1.1666806, 1.1431768, -0.0124158, 2.0594065, 0.1420772, -2.9227523, -2.6610345, -2.0071803, -0.5574015, -1.3192575, -0.8555514, 0.1376866, -2.8049967, -2.2673390, -0.5232039, 1.5473009, -1.2855805, 2.6648289, 1.5906412, 2.5126912, 1.6980225, -2.6334579, 2.8316964, -0.1202799, -2.3108352, -0.7344431, -0.1863690, -0.0075450, 2.9615712, -2.4610171, -0.4309127, -0.4918509, -0.4810587, 2.2077183, -1.4579937, 2.7887593, 2.8904241, -0.1836325, -0.2275295, -0.1299421, 1.2096804, 2.9496770, 1.2184110, 1.2401207, 2.7604226, 0.5534772, -0.0247189, 1.2269684, -2.3566199, -2.9811207, 1.2999521, 0.6409873, -2.7336839, 0.6084908, -2.5626875, 0.5022397, 0.2164019, -2.2245504, 2.1807718, -1.5758820, 2.4466375, 2.0269071, 0.1849097, 2.5777980, -0.5416208, 1.5395423, -0.2795698, -0.5415788, -2.7806202, 2.3278892, -1.5534884, -1.8318555, 0.9536707, -2.2032910, 0.8799313, -1.5041745, -2.3052899, -0.0071255, 1.1934021, -1.9983889, 1.9820110, -1.6687458, 2.7450842, 1.3164705, -2.6535137, 1.2357429, 0.1819178, -1.7003213, -1.6538399, 2.6855732, -0.3064366, 1.7164063, -2.9545294, 2.9010245, -0.0411507, 0.4004713, -2.1868662, 2.5538922, 2.7690421, 2.8188700, -1.7203659, 1.4082227, -1.7725298, -0.1519665, 0.4971974, 2.9286655, -1.3180214, -1.6845799, -2.4987130, 0.0265197, -1.1633564, -1.1011925, 0.1183753, -0.1538756, -1.5842599, -2.7111756, 1.0710594, -2.1830268, 2.6194763, -1.2670836, -1.8177613, -2.7218167, -0.7769317, 2.6260772, 1.9757963, -1.8733269, 2.8810738, -1.6372847, 0.6594904, -2.3871433, -0.2727594, 2.0378350, 2.9517575, 2.8103516, 0.4535808, -2.6226707, -2.2913523, -2.7933397, -0.1644949, -0.9014715, 2.5181358, 1.2539705, -0.7643235, 2.0549231, 2.7802942, -2.8024390, 1.2415348, 0.5538021, -0.8700639, 0.5112655, 0.2984955, -0.3368229, 0.6657549, 0.0070205, -2.1285876, 1.1013324, -1.2674052, -0.1868274, 0.8138506, 2.3955088, -1.1340128, -0.1745562, 0.9361107, 0.3678414, -1.1009564, -2.4152124, -1.7287186, 2.2387078, 1.3284049, 0.1966576, 2.2604411, -0.3887649, 1.2249849, 0.2560314, -1.8728530, 1.4067038, 2.9398708, 0.6421657, 0.7001288, -0.9633487, 2.9304487, 1.4997224, -0.1511689, 0.7525992, -0.3233383, -0.0522308, 0.8805233, 1.1644433, -1.2746032, 0.4484729, 1.8049754, -0.5729506, -1.7219455, -1.3330636, -2.0159999, 0.3768466, -0.1128852, -1.3299456, 0.3609171, -0.1371195, 0.6119481, -2.3379311, 1.8705215, -1.0865461, -1.2860212, -1.5391369, -0.3092695, 1.3184047, 2.1484981, 1.2397678, -1.0321977, 0.6912274, -2.5057045, 1.5010001, -2.3712814, -1.9477828, 0.3249143, 0.5736370, -2.7598556, 2.0707321, -0.6730294, 1.6063768, -1.0398548, 2.3485418, 2.5902571, -2.9208095, 1.6901828, -1.0937468, 1.8212878, -1.8354556, 0.2120741, 2.6987936, -2.1851433, 0.5654253, 1.0269532, -1.4538431, 1.0231416, 2.0811970, -2.4042659, 1.4530665, 1.4192623, -2.1256517, -1.5334988, 0.8556906, 1.4950739, -0.5720348, 0.2919659, 0.2670908, -1.6042114, -1.1645992, -0.7531319, 2.9160717, 0.8665921, -2.3466367, 2.8876809, -0.6324771, -0.6383906, -1.6066410, 1.1110950, 0.9489469, -1.2829955, -2.4665263, 0.8528890, -1.6991289, -0.5491251, 2.7766817, -0.9590528, 1.2870375, 2.5031871, -0.7611168, -1.5965726, -0.5255496, -0.2143821, -1.4976153, 0.2188392, 0.6198784, -0.4349362, 2.4079853, -2.2132712, -0.6589610, 0.8627603, -0.8647738, 0.4696033, -1.6021541, -0.6579570, -1.1940926, -0.6907483, 2.2271030, -2.6160129, -0.6500942, -2.5116133, -1.2402078, 2.1418895, 1.1506459, 0.3916397 );
    constant biases : reals := ( 2.5016475, -0.4769450, -0.4932003, 2.1961096, -2.6706047, 2.3696383, 0.4020859, -1.6265153, -0.3096233, 2.8166511, 1.4735194, 0.1846343, -1.8041594, -2.1763503, -2.9961709, -2.6849192, -2.5794719, 1.4686583, -0.8505542, 2.7954399, 2.1427681, -2.0455065, 0.4455868, 2.0873602, 0.6407637, -2.2499664, 1.9989243, 1.6018489, -0.9843619, -2.3796202, 1.1561464, 2.4479112, -2.5700464, -1.3724784, 2.7492710, 2.9796566, -1.4686636, 2.1163058, 1.5500835, -1.9786676 );
end test_data;
