use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

library work;
use work.util.all;

entity system is
port(
    start : in std_logic;
    test_out : out std_logic_vector(8 - 1 downto 0);
    sel : in unsigned(8 - 1 downto 0)
);
end system;

architecture system of system is

component conv_layer_mc is
generic(
    stride : integer;
    filter_size : integer;
    filter_nb : integer;
    input_size : integer;
    channels : integer;
    dsp_alloc : integer;
    weight_file : string;
    bias_file : string;
    input_int_part : integer;
    input_frac_part : integer;
    weight_int_part : integer;
    weight_frac_part : integer;
    bias_int_part : integer;
    bias_frac_part : integer;
    out_int_part : integer;
    out_frac_part : integer
);
port(
    clk : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    load_done : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    addr : out std_logic_vector;
    out_addr : out std_logic_vector;
    row : out std_logic_vector;
    wren : out std_logic_vector
);
end component;

component bram_pad_interlayer is
generic(
    init_file : string;
    channels : integer;
    channel_width : integer;
    zero_padding : integer;
    layer_size : integer
);
port(
    clk : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    wr_addr : in std_logic_vector;
    rd_addr : in std_logic_vector;
    row : in std_logic_vector;
    wren : in std_logic_vector
);
end component;

component maxpool_layer_mc is
generic(
    pool_size : integer;
    stride : integer;
    input_size : integer;
    channels : integer
);
port(
    clk : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    load_done : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    addr : out std_logic_vector;
    out_addr : out std_logic_vector;
    row : out std_logic_vector;
    wren : out std_logic_vector
);
end component;

component fc_layer is
generic(
    input_width : integer;
    output_width : integer;
    simd_width : integer;
    input_spec : fixed_spec;
    weight_spec : fixed_spec;
    op_arg_spec : fixed_spec;
    output_spec : fixed_spec;
    n_weights : integer;
    pick_from_ram : boolean;
    weights_filename : string;
    weight_values : reals
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    in_a : in std_logic_vector;
    out_a : out std_logic_vector;
    out_offset : out unsigned;
    simd_offset : out std_logic_vector;
    op_argument : out sfixed;
    op_result : in sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component conv_to_fc_interlayer is
generic(
    channels : integer;
    channel_width : integer;
    layer_size : integer;
    fc_simd : integer
);
port(
    clk : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    ack : out std_logic;
    din : in std_logic_vector;
    dout : out std_logic_vector;
    wr_addr : in std_logic_vector;
    rd_addr : in std_logic_vector;
    wren_in : in std_logic_vector
);
end component;

component bias_op is
generic(
    input_spec : fixed_spec;
    bias_spec : fixed_spec;
    biases : reals
);
port(
    input : in sfixed;
    offset : in unsigned;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component sigmoid_op is
generic(
    input_spec : fixed_spec;
    output_spec : fixed_spec;
    step_precision : integer;
    bit_precision : integer
);
port(
    clk : in std_logic;
    input : in sfixed;
    output : out sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;



signal ready_s1 : std_logic;
signal done_s2 : std_logic;
signal start_s3 : std_logic;
signal ack_s4 : std_logic;
signal load_done_s5 : std_logic;
signal din_s6 : std_logic_vector(7 downto 0);
signal dout_s7 : std_logic_vector(79 downto 0);
signal addr_s8 : std_logic_vector(9 downto 0);
signal out_addr_s9 : std_logic_vector(9 downto 0);
signal row_s10 : std_logic_vector(4 downto 0);
signal wren_s11 : std_logic_vector(9 downto 0);


signal ready_s74 : std_logic;
signal done_s75 : std_logic;
signal start_s76 : std_logic;
signal din_s77 : std_logic_vector(7 downto 0);
signal dout_s78 : std_logic_vector(7 downto 0);
signal wr_addr_s79 : std_logic_vector(9 downto 0);
signal rd_addr_s80 : std_logic_vector(9 downto 0);
signal row_s81 : std_logic_vector(4 downto 0);
signal wren_s82 : std_logic_vector(0 downto 0);


signal ready_s13 : std_logic;
signal done_s14 : std_logic;
signal start_s15 : std_logic;
signal ack_s16 : std_logic;
signal load_done_s17 : std_logic;
signal din_s18 : std_logic_vector(79 downto 0);
signal dout_s19 : std_logic_vector(79 downto 0);
signal addr_s20 : std_logic_vector(9 downto 0);
signal out_addr_s21 : std_logic_vector(7 downto 0);
signal row_s22 : std_logic_vector(3 downto 0);
signal wren_s23 : std_logic_vector(9 downto 0);


signal ready_s84 : std_logic;
signal done_s85 : std_logic;
signal start_s86 : std_logic;
signal din_s87 : std_logic_vector(79 downto 0);
signal dout_s88 : std_logic_vector(79 downto 0);
signal wr_addr_s89 : std_logic_vector(9 downto 0);
signal rd_addr_s90 : std_logic_vector(9 downto 0);
signal row_s91 : std_logic_vector(4 downto 0);
signal wren_s92 : std_logic_vector(9 downto 0);


signal ready_s25 : std_logic;
signal done_s26 : std_logic;
signal start_s27 : std_logic;
signal ack_s28 : std_logic;
signal load_done_s29 : std_logic;
signal din_s30 : std_logic_vector(79 downto 0);
signal dout_s31 : std_logic_vector(79 downto 0);
signal addr_s32 : std_logic_vector(8 downto 0);
signal out_addr_s33 : std_logic_vector(7 downto 0);
signal row_s34 : std_logic_vector(3 downto 0);
signal wren_s35 : std_logic_vector(9 downto 0);


signal ready_s94 : std_logic;
signal done_s95 : std_logic;
signal start_s96 : std_logic;
signal din_s97 : std_logic_vector(79 downto 0);
signal dout_s98 : std_logic_vector(79 downto 0);
signal wr_addr_s99 : std_logic_vector(7 downto 0);
signal rd_addr_s100 : std_logic_vector(8 downto 0);
signal row_s101 : std_logic_vector(3 downto 0);
signal wren_s102 : std_logic_vector(9 downto 0);


signal ready_s37 : std_logic;
signal done_s38 : std_logic;
signal start_s39 : std_logic;
signal ack_s40 : std_logic;
signal load_done_s41 : std_logic;
signal din_s42 : std_logic_vector(79 downto 0);
signal dout_s43 : std_logic_vector(79 downto 0);
signal addr_s44 : std_logic_vector(7 downto 0);
signal out_addr_s45 : std_logic_vector(5 downto 0);
signal row_s46 : std_logic_vector(2 downto 0);
signal wren_s47 : std_logic_vector(9 downto 0);


signal ready_s104 : std_logic;
signal done_s105 : std_logic;
signal start_s106 : std_logic;
signal din_s107 : std_logic_vector(79 downto 0);
signal dout_s108 : std_logic_vector(79 downto 0);
signal wr_addr_s109 : std_logic_vector(7 downto 0);
signal rd_addr_s110 : std_logic_vector(7 downto 0);
signal row_s111 : std_logic_vector(3 downto 0);
signal wren_s112 : std_logic_vector(9 downto 0);



signal ready_s49 : std_logic;
signal done_s50 : std_logic;
signal start_s51 : std_logic;
signal ack_s52 : std_logic;
signal in_a_s53 : std_logic_vector(89 downto 0);
signal out_a_s54 : std_logic_vector(99 downto 0);
signal out_offset_s55 : unsigned(3 downto 0);
signal simd_offset_s56 : std_logic_vector(5 downto 0);
signal op_argument_s57 : sfixed(12 downto -15);
signal op_result_s58 : sfixed(1 downto -8);
signal op_send_s59 : std_logic;
signal op_receive_s60 : std_logic;


signal ready_s115 : std_logic;
signal done_s116 : std_logic;
signal start_s117 : std_logic;
signal ack_s118 : std_logic;
signal din_s119 : std_logic_vector(79 downto 0);
signal dout_s120 : std_logic_vector(89 downto 0);
signal wr_addr_s121 : std_logic_vector(5 downto 0);
signal rd_addr_s122 : std_logic_vector(0 downto 0);
signal wren_in_s123 : std_logic_vector(9 downto 0);

signal input_s62 : sfixed(12 downto -15);
signal offset_s63 : unsigned(3 downto 0);
signal output_s64 : sfixed(13 downto -15);
signal op_send_s65 : std_logic;
signal op_receive_s66 : std_logic;


signal input_s68 : sfixed(13 downto -15);
signal output_s69 : sfixed(1 downto -8);
signal op_send_s70 : std_logic;
signal op_receive_s71 : std_logic;


component ps_clk is
port(
    clk, rst : out std_logic
);
end component;

signal clk, rst_sink : std_logic;
constant rst : std_logic := '0';


begin

conv_layer_mc_u0 : conv_layer_mc generic map(
    stride => 1,
    filter_size => 5,
    filter_nb => 10,
    input_size => 32,
    channels => 1,
    dsp_alloc => 1,
    weight_file => "C:/Users/gademb/stage2017/Gabriel/codegen/convgentest/conv-w1.nn",
    bias_file => "C:/Users/gademb/stage2017/Gabriel/codegen/convgentest/conv-b1.nn",
    input_int_part => 0,
    input_frac_part => 8,
    weight_int_part => 1,
    weight_frac_part => 8,
    bias_int_part => 1,
    bias_frac_part => 8,
    out_int_part => 0,
    out_frac_part => 8
) port map(
    clk => clk,
    ready => ready_s1,
    done => done_s2,
    start => start_s3,
    ack => ack_s4,
    load_done => load_done_s5,
    din => din_s6,
    dout => dout_s7,
    addr => addr_s8,
    out_addr => out_addr_s9,
    row => row_s10,
    wren => wren_s11
);
bram_pad_interlayer_u73 : bram_pad_interlayer generic map(
    init_file => "C:/Users/gademb/stage2017/Gabriel/codegen/convgentest/conv-b1.nn",
    channels => 1,
    channel_width => 8,
    zero_padding => 2,
    layer_size => 28
) port map(
    clk => clk,
    ready => ready_s74,
    done => done_s75,
    start => start_s76,
    din => din_s77,
    dout => dout_s78,
    wr_addr => wr_addr_s79,
    rd_addr => rd_addr_s80,
    row => row_s81,
    wren => wren_s82
);
maxpool_layer_mc_u12 : maxpool_layer_mc generic map(
    pool_size => 2,
    stride => 2,
    input_size => 28,
    channels => 10
) port map(
    clk => clk,
    ready => ready_s13,
    done => done_s14,
    start => start_s15,
    ack => ack_s16,
    load_done => load_done_s17,
    din => din_s18,
    dout => dout_s19,
    addr => addr_s20,
    out_addr => out_addr_s21,
    row => row_s22,
    wren => wren_s23
);
bram_pad_interlayer_u83 : bram_pad_interlayer generic map(
    init_file => "",
    channels => 10,
    channel_width => 8,
    zero_padding => 0,
    layer_size => 28
) port map(
    clk => clk,
    ready => ready_s84,
    done => done_s85,
    start => start_s86,
    din => din_s87,
    dout => dout_s88,
    wr_addr => wr_addr_s89,
    rd_addr => rd_addr_s90,
    row => row_s91,
    wren => wren_s92
);
conv_layer_mc_u24 : conv_layer_mc generic map(
    stride => 1,
    filter_size => 5,
    filter_nb => 10,
    input_size => 18,
    channels => 10,
    dsp_alloc => 5,
    weight_file => "C:/Users/gademb/stage2017/Gabriel/codegen/convgentest/conv-w2.nn",
    bias_file => "C:/Users/gademb/stage2017/Gabriel/codegen/convgentest/conv-b2.nn",
    input_int_part => 0,
    input_frac_part => 8,
    weight_int_part => 1,
    weight_frac_part => 8,
    bias_int_part => 1,
    bias_frac_part => 8,
    out_int_part => 0,
    out_frac_part => 8
) port map(
    clk => clk,
    ready => ready_s25,
    done => done_s26,
    start => start_s27,
    ack => ack_s28,
    load_done => load_done_s29,
    din => din_s30,
    dout => dout_s31,
    addr => addr_s32,
    out_addr => out_addr_s33,
    row => row_s34,
    wren => wren_s35
);
bram_pad_interlayer_u93 : bram_pad_interlayer generic map(
    init_file => "",
    channels => 10,
    channel_width => 8,
    zero_padding => 2,
    layer_size => 14
) port map(
    clk => clk,
    ready => ready_s94,
    done => done_s95,
    start => start_s96,
    din => din_s97,
    dout => dout_s98,
    wr_addr => wr_addr_s99,
    rd_addr => rd_addr_s100,
    row => row_s101,
    wren => wren_s102
);
maxpool_layer_mc_u36 : maxpool_layer_mc generic map(
    pool_size => 2,
    stride => 2,
    input_size => 14,
    channels => 10
) port map(
    clk => clk,
    ready => ready_s37,
    done => done_s38,
    start => start_s39,
    ack => ack_s40,
    load_done => load_done_s41,
    din => din_s42,
    dout => dout_s43,
    addr => addr_s44,
    out_addr => out_addr_s45,
    row => row_s46,
    wren => wren_s47
);
bram_pad_interlayer_u103 : bram_pad_interlayer generic map(
    init_file => "",
    channels => 10,
    channel_width => 8,
    zero_padding => 0,
    layer_size => 14
) port map(
    clk => clk,
    ready => ready_s104,
    done => done_s105,
    start => start_s106,
    din => din_s107,
    dout => dout_s108,
    wr_addr => wr_addr_s109,
    rd_addr => rd_addr_s110,
    row => row_s111,
    wren => wren_s112
);
fc_layer_u48 : fc_layer generic map(
    input_width => 490,
    output_width => 10,
    simd_width => 10,
    input_spec => fixed_spec(fixed_spec'(int => 1, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 1, frac => 7)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 13, frac => 15)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    n_weights => 31360,
    pick_from_ram => true,
    weights_filename => "whatever",
    weight_values => reals(reals'( 0.2580850, 0.6637810, 0.7317050, 0.9346510, 0.5235030, 0.3026220, 0.6658780, 0.1178690, 0.3872960, 0.7304440, 0.1125770, 0.1015950, 0.5039400, 0.1663390, 0.7121680, 0.3713270, 0.8353030, 0.6779000, 0.0287057, 0.8338360, 0.3615540, 0.3427120, 0.5462880, 0.6234020, 0.0226888, 0.5343000, 0.1493000, 0.5142030, 0.6155320, 0.0931069, 0.4533790, 0.6693380, 0.5207680, 0.9990630, 0.0484407, 0.7212360, 0.8510440, 0.9121590, 0.6477040, 0.9708820, 0.9900710, 0.5097420, 0.1019290, 0.6708780, 0.9406110, 0.2308030, 0.9592590, 0.7907010, 0.0907339, 0.7214400, 0.5751610, 0.9607440, 0.0466014, 0.7676290, 0.3457780, 0.7744330, 0.2014980, 0.8479960, 0.5127080, 0.6629040, 0.5919950, 0.5667360, 0.7718270, 0.2223950, 0.1956730, 0.7298820, 0.9010540, 0.0271075, 0.0706680, 0.8253170, 0.8854490, 0.1468050, 0.3334790, 0.0198137, 0.1212620, 0.0554147, 0.6474440, 0.5228840, 0.9029290, 0.7045460, 0.3488960, 0.1924570, 0.6426200, 0.7189440, 0.4708310, 0.7257350, 0.0012637, 0.5738260, 0.9783650, 0.5077320, 0.8764130, 0.2144910, 0.0202081, 0.6061750, 0.5166570, 0.9961360, 0.6846190, 0.0017873, 0.0556836, 0.7787720, 0.2356630, 0.9033550, 0.6182470, 0.8203120, 0.8496210, 0.6960010, 0.4944680, 0.0014134, 0.6543350, 0.4190760, 0.1537620, 0.2684350, 0.5233300, 0.1164910, 0.1498260, 0.6478090, 0.2413950, 0.6246050, 0.3734960, 0.1306520, 0.0137214, 0.0785052, 0.3579070, 0.3902330, 0.8740390, 0.7819720, 0.1787390, 0.1388680, 0.9094710, 0.5438470, 0.6315710, 0.2811350, 0.1999680, 0.4450670, 0.0096940, 0.8370290, 0.2733950, 0.8099340, 0.8529010, 0.1801690, 0.3020440, 0.0505371, 0.8588310, 0.3175110, 0.7636410, 0.7984670, 0.8225900, 0.0154416, 0.7075900, 0.0875132, 0.7831210, 0.4934420, 0.1431200, 0.8459540, 0.7790000, 0.4824980, 0.7974080, 0.3039870, 0.4116160, 0.1819620, 0.8188600, 0.9903160, 0.0272449, 0.4357500, 0.7893190, 0.3904540, 0.4099020, 0.0471540, 0.5120500, 0.3340420, 0.7280580, 0.4102690, 0.3640820, 0.8335600, 0.6997870, 0.7196660, 0.4357960, 0.0095928, 0.6290550, 0.2776610, 0.6976570, 0.0166568, 0.8626900, 0.4646260, 0.6207130, 0.3555190, 0.5558570, 0.4253690, 0.7034130, 0.9616890, 0.9326640, 0.1218820, 0.4742730, 0.7924200, 0.9000000, 0.7695290, 0.3779270, 0.2429200, 0.5016840, 0.3336460, 0.7986230, 0.5145470, 0.8708940, 0.7334320, 0.4095870, 0.1764820, 0.7656470, 0.9592760, 0.2166980, 0.9962180, 0.0875456, 0.8488650, 0.1683630, 0.6863830, 0.8784540, 0.7687470, 0.8353720, 0.5044110, 0.3463660, 0.8248240, 0.6352960, 0.8888660, 0.6202730, 0.8772590, 0.7513180, 0.5949840, 0.2300010, 0.8896740, 0.3219950, 0.9499280, 0.8578010, 0.8167540, 0.4879290, 0.9207930, 0.8048020, 0.9919180, 0.3460190, 0.8740890, 0.4520540, 0.9327930, 0.1884010, 0.1462720, 0.0699236, 0.1849910, 0.0396100, 0.1500420, 0.1142610, 0.4974280, 0.5631420, 0.8776930, 0.4500250, 0.5913660, 0.9119600, 0.4775020, 0.0733154, 0.4576770, 0.1594620, 0.9082380, 0.0235826, 0.9495190, 0.7762930, 0.3373530, 0.6337600, 0.1496760, 0.2077700, 0.7005190, 0.0396725, 0.4181710, 0.7681340, 0.3537960, 0.3430990, 0.8178110, 0.8506070, 0.6781000, 0.5882190, 0.0407057, 0.7228330, 0.8629690, 0.5145510, 0.9028630, 0.7733110, 0.1575680, 0.4726600, 0.0740094, 0.9688150, 0.7500560, 0.7156540, 0.4469810, 0.9739810, 0.2271300, 0.0279454, 0.4559110, 0.3846820, 0.5889000, 0.1160140, 0.0976037, 0.4474040, 0.7457900, 0.4103040, 0.0076341, 0.9958870, 0.6159550, 0.5262110, 0.2873580, 0.8814220, 0.2585070, 0.1174600, 0.1041670, 0.7213340, 0.9819890, 0.3164110, 0.1193480, 0.4717360, 0.7688670, 0.5847000, 0.2488700, 0.4210150, 0.2399100, 0.0063004, 0.0065578, 0.8079270, 0.1187150, 0.3880040, 0.1072320, 0.7302490, 0.4130320, 0.9140080, 0.4652290, 0.1579550, 0.2776600, 0.8328600, 0.6528290, 0.8649970, 0.9129140, 0.4276910, 0.2041230, 0.5245470, 0.5454110, 0.7671390, 0.0973710, 0.9166420, 0.0578557, 0.6428590, 0.5486520, 0.7557970, 0.1313700, 0.9702860, 0.1452980, 0.5674660, 0.1230020, 0.7102310, 0.1990510, 0.4103760, 0.4546310, 0.6704910, 0.7420830, 0.0507930, 0.2704100, 0.5881900, 0.6931590, 0.9973310, 0.5056820, 0.1166410, 0.7125960, 0.4933250, 0.4271240, 0.7274010, 0.7761610, 0.2847950, 0.0525871, 0.5882310, 0.0005306, 0.7242180, 0.6208550, 0.4475710, 0.0056616, 0.3679100, 0.1640770, 0.8279710, 0.6407940, 0.2916390, 0.8771380, 0.6345140, 0.2038980, 0.1481480, 0.8181930, 0.2987750, 0.2459800, 0.0823575, 0.9830570, 0.1476230, 0.8886480, 0.5397910, 0.4519430, 0.0042354, 0.9361250, 0.2745860, 0.7466700, 0.0742473, 0.2882950, 0.6181650, 0.5161480, 0.3176020, 0.4532280, 0.4648930, 0.5818200, 0.8156290, 0.8946450, 0.9761350, 0.9679390, 0.1254660, 0.2304830, 0.7883160, 0.8322780, 0.3954860, 0.7299650, 0.5720020, 0.5384660, 0.3749090, 0.1873650, 0.2888640, 0.0318466, 0.8041680, 0.7191960, 0.4977020, 0.2596010, 0.1338940, 0.2649130, 0.8162770, 0.6901240, 0.3912210, 0.7359440, 0.7069400, 0.1788960, 0.5290830, 0.0794923, 0.1386910, 0.5696120, 0.9239490, 0.3120910, 0.9724780, 0.9023800, 0.6701370, 0.0228402, 0.3820770, 0.1628390, 0.5057150, 0.5467200, 0.6655350, 0.4604970, 0.8027720, 0.0994835, 0.0996270, 0.8589120, 0.1123310, 0.6290670, 0.5051840, 0.5622840, 0.2163750, 0.0614157, 0.8424270, 0.6730270, 0.4872010, 0.3423820, 0.5286200, 0.6194170, 0.3301720, 0.2364320, 0.4985810, 0.1387260, 0.5630870, 0.1617270, 0.0150216, 0.3403820, 0.4017540, 0.5350040, 0.0919819, 0.1251600, 0.7339700, 0.5321960, 0.7031020, 0.0794658, 0.1308030, 0.9901450, 0.3842820, 0.2908490, 0.8344040, 0.6876760, 0.0807336, 0.9798110, 0.5385450, 0.2215850, 0.8062640, 0.0230655, 0.8999200, 0.7756830, 0.6468900, 0.6535220, 0.8201370, 0.4928370, 0.3812430, 0.9058800, 0.9091710, 0.9642920, 0.3727960, 0.6359920, 0.3592800, 0.2999390, 0.4126640, 0.3483440, 0.0309225, 0.3828580, 0.3791910, 0.0345070, 0.4366330, 0.8066700, 0.3029050, 0.8304280, 0.9123080, 0.4909290, 0.3021190, 0.2368390, 0.6841430, 0.0367383, 0.2153850, 0.9863770, 0.9513140, 0.5682800, 0.6779910, 0.9771710, 0.7305070, 0.4203440, 0.7020000, 0.8321630, 0.0775366, 0.1253610, 0.4454040, 0.3569910, 0.1442000, 0.9120100, 0.6092890, 0.3925250, 0.9580570, 0.8670750, 0.6798080, 0.3046870, 0.7570160, 0.7946360, 0.6749110, 0.8335150, 0.6505330, 0.2276160, 0.5005670, 0.7948330, 0.4865140, 0.5792580, 0.2207050, 0.4000320, 0.4198420, 0.5230640, 0.9799970, 0.8556760, 0.0884017, 0.9990910, 0.7708070, 0.1364670, 0.7012510, 0.7245980, 0.1423630, 0.0551354, 0.1263970, 0.7362760, 0.1675820, 0.7909280, 0.5743120, 0.5820780, 0.2536130, 0.6126470, 0.1948400, 0.4357240, 0.0987317, 0.8848750, 0.9830360, 0.5171040, 0.6141710, 0.6406660, 0.3293240, 0.1219240, 0.1309850, 0.3420820, 0.9309030, 0.4457170, 0.9091250, 0.7088070, 0.1743870, 0.3796770, 0.3762410, 0.5012560, 0.8147170, 0.7158630, 0.9235460, 0.0004639, 0.3914120, 0.0494234, 0.5295920, 0.8890700, 0.5794020, 0.2265150, 0.6668230, 0.8271820, 0.2345940, 0.7623510, 0.0001186, 0.5320480, 0.4083620, 0.7716890, 0.2365970, 0.9823090, 0.2139040, 0.0392147, 0.4624910, 0.5463810, 0.4390150, 0.7092100, 0.1983350, 0.7640130, 0.1455990, 0.6137700, 0.1397680, 0.3869840, 0.3897600, 0.6237600, 0.8031110, 0.6618720, 0.7095480, 0.1926630, 0.0692082, 0.5975890, 0.4170450, 0.7533010, 0.2928190, 0.3063900, 0.1777050, 0.9892490, 0.6535230, 0.5679220, 0.0163062, 0.6648690, 0.5729990, 0.2752330, 0.8587300, 0.9534870, 0.5028880, 0.1967370, 0.8917090, 0.1478370, 0.4957080, 0.2192370, 0.4934360, 0.7856620, 0.8756370, 0.3243670, 0.4019580, 0.7203340, 0.1797170, 0.8895330, 0.3926510, 0.9317360, 0.7398150, 0.2469540, 0.0666942, 0.4572340, 0.7158300, 0.9199360, 0.4819890, 0.4361840, 0.3214410, 0.7827470, 0.5709070, 0.2327980, 0.9366780, 0.1258060, 0.5292700, 0.2834000, 0.6024990, 0.2565480, 0.7276560, 0.9287360, 0.1255440, 0.9868320, 0.6228390, 0.6577870, 0.7055830, 0.8392860, 0.9533680, 0.6041760, 0.7003170, 0.8738560, 0.3614020, 0.8469690, 0.4600440, 0.7390880, 0.2975370, 0.2588520, 0.2127660, 0.6147130, 0.1966000, 0.2590260, 0.5429540, 0.9520540, 0.4385280, 0.4046250, 0.0427279, 0.0478010, 0.0892147, 0.4345650, 0.7893120, 0.1931000, 0.8231960, 0.4886040, 0.7840420, 0.2913260, 0.1277000, 0.6718080, 0.0125924, 0.1159200, 0.0082810, 0.3929610, 0.0892128, 0.9200390, 0.6832620, 0.8976210, 0.4700120, 0.4486960, 0.4942670, 0.9111750, 0.5948060, 0.1283570, 0.7688900, 0.5015110, 0.8494270, 0.2570830, 0.3660330, 0.5081220, 0.9850780, 0.6725720, 0.2937900, 0.1704090, 0.0977367, 0.0626736, 0.8694380, 0.7848980, 0.4538710, 0.5987540, 0.9205860, 0.7427720, 0.5264070, 0.9302990, 0.3937770, 0.1957580, 0.6559040, 0.3880360, 0.3173840, 0.2680780, 0.0935761, 0.2895330, 0.6215810, 0.4465090, 0.4051700, 0.5383740, 0.4206640, 0.1756460, 0.4242160, 0.2608800, 0.9597060, 0.5458150, 0.0359280, 0.7770410, 0.4124920, 0.9389960, 0.2987840, 0.7100560, 0.8366910, 0.1380430, 0.2227290, 0.3379350, 0.0952702, 0.6139090, 0.6423190, 0.3191600, 0.5185120, 0.4736900, 0.7366330, 0.6680290, 0.6379640, 0.5972150, 0.8001400, 0.5839980, 0.1129000, 0.1421650, 0.7225410, 0.0981930, 0.9629310, 0.8830920, 0.2735620, 0.1747210, 0.2933380, 0.7897320, 0.7685620, 0.9766190, 0.3152760, 0.6483520, 0.7655060, 0.5858170, 0.5191190, 0.0921713, 0.0828014, 0.9455480, 0.1129090, 0.1069580, 0.1196150, 0.8171490, 0.7747240, 0.7422520, 0.5115140, 0.4717080, 0.4736690, 0.5521190, 0.4262130, 0.7142430, 0.7416640, 0.1466000, 0.0777698, 0.8176730, 0.2056190, 0.6365130, 0.1588290, 0.2893960, 0.7272990, 0.2178290, 0.0521419, 0.9145820, 0.7701840, 0.0248357, 0.1066610, 0.6471670, 0.4748980, 0.2002310, 0.3613170, 0.6933590, 0.1831560, 0.4084630, 0.3054920, 0.6014740, 0.3362210, 0.8747420, 0.7918380, 0.1635010, 0.0870523, 0.2163950, 0.0285462, 0.9481400, 0.1189500, 0.9876190, 0.4447770, 0.6183110, 0.5152310, 0.6073100, 0.1271600, 0.7002060, 0.2006620, 0.0438648, 0.6918390, 0.3623210, 0.4232640, 0.9329690, 0.3017100, 0.2468420, 0.2454880, 0.9177600, 0.5914140, 0.2725680, 0.6289130, 0.5972070, 0.2336790, 0.9844680, 0.5438750, 0.6518350, 0.5256580, 0.3766590, 0.1895930, 0.5715490, 0.9613530, 0.6559750, 0.9588190, 0.4293660, 0.0745202, 0.5028590, 0.6530170, 0.6088960, 0.6799220, 0.4388330, 0.0815753, 0.0325830, 0.1204070, 0.2679180, 0.7259720, 0.9394950, 0.6870350, 0.7090660, 0.5418140, 0.4914540, 0.2320530, 0.9824810, 0.3508830, 0.0018719, 0.7920730, 0.4943910, 0.1017250, 0.4279690, 0.8040370, 0.6877520, 0.5991220, 0.9341370, 0.7593610, 0.2561840, 0.3041270, 0.0823527, 0.9189170, 0.1851200, 0.1421220, 0.1044750, 0.8388480, 0.1085950, 0.0259800, 0.6709430, 0.6632400, 0.7397110, 0.7711070, 0.1893740, 0.2631810, 0.8767720, 0.7579410, 0.9872690, 0.4538440, 0.2285140, 0.0791225, 0.4160330, 0.1552400, 0.7075390, 0.0502966, 0.3523970, 0.2462010, 0.1406120, 0.6703580, 0.0042149, 0.0075302, 0.7612600, 0.7040720, 0.0399742, 0.1477850, 0.2272190, 0.3332590, 0.7991860, 0.6878760, 0.3440980, 0.5920150, 0.7525020, 0.9944850, 0.3891330, 0.0965254, 0.6369670, 0.1856310, 0.5587860, 0.2344930, 0.7190570, 0.5957970, 0.0602838, 0.1629980, 0.3556870, 0.0871918, 0.4980470, 0.9960120, 0.3246300, 0.8241510, 0.3173870, 0.9920680, 0.2748230, 0.3282770, 0.3295200, 0.2224420, 0.0524683, 0.9822530, 0.6678730, 0.8010320, 0.6590520, 0.2318010, 0.9327050, 0.1396580, 0.9498150, 0.9646420, 0.1815190, 0.3759630, 0.5191730, 0.9302510, 0.2030540, 0.2291650, 0.0479666, 0.2115820, 0.2713800, 0.8490010, 0.6822570, 0.5184810, 0.5458860, 0.1752400, 0.2967630, 0.1886870, 0.6660590, 0.7168560, 0.2090080, 0.7201050, 0.1235770, 0.9751690, 0.3520250, 0.0205234, 0.9560510, 0.6878840, 0.0583234, 0.9287740, 0.0622763, 0.2574730, 0.0652294, 0.9321560, 0.3982220, 0.4240920, 0.3170560, 0.3855070, 0.7978050, 0.7835780, 0.7887360, 0.9914210, 0.7288420, 0.4856920, 0.1793390, 0.8685180, 0.6264050, 0.7824860, 0.7270890, 0.1922810, 0.0001228, 0.0333845, 0.2257350, 0.8814130, 0.6110990, 0.6884240, 0.4702800, 0.6466980, 0.5555200, 0.7627460, 0.2462270, 0.1857880, 0.4035730, 0.7523120, 0.0192597, 0.7398250, 0.7863510, 0.6530320, 0.0695931, 0.2255790, 0.8218940, 0.4113130, 0.7619200, 0.0857349, 0.7288680, 0.8311210, 0.2535750, 0.7340390, 0.7573110, 0.5033270, 0.9086360, 0.0575505, 0.4174280, 0.6508500, 0.7759280, 0.8664520, 0.8885530, 0.1704100, 0.0635901, 0.3143530, 0.8694690, 0.5085470, 0.7289810, 0.5255370, 0.1605590, 0.8352700, 0.9655360, 0.4679920, 0.7445780, 0.2580560, 0.3444330, 0.5394620, 0.0184294, 0.8126450, 0.6041130, 0.4483720, 0.4313700, 0.8857160, 0.9775940, 0.5153750, 0.1514020, 0.5054720, 0.4459830, 0.6319370, 0.4177580, 0.6678390, 0.4632790, 0.5409370, 0.1754710, 0.4436950, 0.8366100, 0.7300140, 0.6665500, 0.4851460, 0.1372350, 0.1501140, 0.4692520, 0.8999820, 0.7346150, 0.4096160, 0.2215760, 0.0786305, 0.6635910, 0.4511260, 0.1880500, 0.0124545, 0.1689350, 0.6494340, 0.6813490, 0.6384990, 0.6803160, 0.1847340, 0.3566890, 0.0879301, 0.7192940, 0.5783770, 0.9164850, 0.9175020, 0.5107250, 0.5782780, 0.8069550, 0.8629750, 0.5286230, 0.5060570, 0.4074430, 0.6504990, 0.6370850, 0.5522620, 0.1722990, 0.7897650, 0.5670970, 0.6842220, 0.3894910, 0.7013380, 0.9056870, 0.6036730, 0.6366630, 0.3313210, 0.4081720, 0.8639740, 0.8006110, 0.1063080, 0.8288660, 0.2505710, 0.1550460, 0.6534620, 0.1892980, 0.1776290, 0.0231114, 0.4731170, 0.3394940, 0.3390360, 0.7586390, 0.4220240, 0.7344260, 0.8126050, 0.5682770, 0.3585830, 0.4427690, 0.3130740, 0.4296670, 0.6188620, 0.1944110, 0.4053430, 0.7171130, 0.6385480, 0.2606050, 0.8910040, 0.1058150, 0.4992100, 0.4708630, 0.5436340, 0.2578990, 0.8250370, 0.1403860, 0.3277250, 0.9460990, 0.9953280, 0.6384700, 0.7844740, 0.1814870, 0.8028190, 0.4345190, 0.7007560, 0.4829670, 0.8465000, 0.1623500, 0.3442380, 0.9707450, 0.0254355, 0.2926190, 0.1112920, 0.4673620, 0.0092502, 0.9722610, 0.6420550, 0.3759330, 0.9440810, 0.2320860, 0.1522730, 0.5897810, 0.3264210, 0.8160530, 0.0548715, 0.0147836, 0.4589690, 0.0472404, 0.2656210, 0.8133550, 0.6503520, 0.4140620, 0.6782570, 0.3200800, 0.5182870, 0.3347390, 0.5839270, 0.1272770, 0.4652510, 0.0310846, 0.3087760, 0.4015710, 0.8054530, 0.2767860, 0.2283010, 0.5384700, 0.3426470, 0.6536890, 0.3722970, 0.8512600, 0.3418010, 0.6191510, 0.3481930, 0.2487180, 0.6037900, 0.2797030, 0.6534160, 0.3029090, 0.3862900, 0.9206890, 0.4169860, 0.6810590, 0.2982380, 0.2604260, 0.6502260, 0.8464720, 0.7860600, 0.2438590, 0.4728060, 0.2691710, 0.0753054, 0.2011340, 0.1477220, 0.7154420, 0.6871750, 0.0464744, 0.6417580, 0.5828440, 0.8291510, 0.0079106, 0.3253290, 0.9683380, 0.8783340, 0.0925172, 0.4753590, 0.4768400, 0.6215420, 0.3406490, 0.0843924, 0.6845030, 0.8401080, 0.9528870, 0.1575160, 0.4482510, 0.2606040, 0.8877150, 0.9260440, 0.3687730, 0.1291290, 0.4425770, 0.0976070, 0.8843730, 0.4893400, 0.7530160, 0.9818690, 0.5403220, 0.3944340, 0.5024650, 0.2129850, 0.1989550, 0.3878310, 0.0319314, 0.6916170, 0.4318810, 0.1786300, 0.7615490, 0.1739340, 0.1057650, 0.7961110, 0.8148960, 0.7393590, 0.7891880, 0.4743410, 0.1030150, 0.8360830, 0.9149840, 0.3794970, 0.8474800, 0.8428390, 0.7144100, 0.8076620, 0.7585230, 0.3363530, 0.7445300, 0.8044720, 0.7785020, 0.6936500, 0.9890660, 0.5892360, 0.9433090, 0.9248070, 0.8563060, 0.1143950, 0.3287530, 0.2995840, 0.5071900, 0.2836830, 0.8448720, 0.1567510, 0.8284880, 0.9380470, 0.5591160, 0.2621800, 0.4946380, 0.6284710, 0.2302850, 0.3303330, 0.5183740, 0.8864970, 0.7396070, 0.8927480, 0.0393736, 0.8965910, 0.5715860, 0.8164240, 0.3851560, 0.4022310, 0.5280840, 0.5433610, 0.8247310, 0.0598475, 0.8524320, 0.6073050, 0.2117360, 0.8800320, 0.3090050, 0.8492660, 0.3560130, 0.0541623, 0.8496670, 0.5828130, 0.5137830, 0.8223350, 0.8976790, 0.2665180, 0.9143360, 0.9859140, 0.4039500, 0.2090320, 0.7817920, 0.2679180, 0.2961850, 0.4228860, 0.0474241, 0.0423018, 0.4635640, 0.0498388, 0.7622430, 0.7970580, 0.2172340, 0.8417130, 0.7306790, 0.0032494, 0.3458990, 0.7417240, 0.2050030, 0.3272690, 0.9795930, 0.9573710, 0.2263250, 0.5472660, 0.7835200, 0.6472560, 0.4681740, 0.0796530, 0.7524810, 0.9512460, 0.7119320, 0.7357030, 0.8333530, 0.0052110, 0.2786360, 0.3406900, 0.0909812, 0.8495850, 0.0439774, 0.4706950, 0.9460340, 0.5166490, 0.4702160, 0.1495720, 0.3155860, 0.1038920, 0.1353220, 0.8412770, 0.0559217, 0.7218220, 0.1664500, 0.0452311, 0.4735560, 0.9121560, 0.6077700, 0.1597120, 0.2220350, 0.9759830, 0.9641870, 0.1876070, 0.9402130, 0.7285770, 0.9164450, 0.0160764, 0.2794150, 0.8961660, 0.2302630, 0.7354120, 0.1148630, 0.7289440, 0.7738650, 0.6891710, 0.1970290, 0.4537940, 0.2906790, 0.3714520, 0.8777910, 0.0205314, 0.6310060, 0.8365250, 0.9563440, 0.3974640, 0.2506010, 0.8107380, 0.1408620, 0.9067570, 0.1908860, 0.0714416, 0.4558740, 0.9611190, 0.9449840, 0.2784000, 0.6683330, 0.8653150, 0.2464340, 0.3584710, 0.3492060, 0.7046840, 0.3013900, 0.8936290, 0.2751470, 0.7036190, 0.8702200, 0.1477400, 0.9809730, 0.2202800, 0.4655900, 0.6600380, 0.2935580, 0.0960612, 0.7015270, 0.0475337, 0.9527930, 0.4850660, 0.1317790, 0.3145040, 0.8059240, 0.4934260, 0.3269360, 0.8549670, 0.3605010, 0.3144030, 0.4630120, 0.0775238, 0.3189140, 0.4503710, 0.1118790, 0.2385110, 0.3140520, 0.0435392, 0.6611690, 0.3013520, 0.1889740, 0.8760970, 0.3766820, 0.1400160, 0.3091530, 0.3302190, 0.6657830, 0.3415880, 0.7481160, 0.4704370, 0.9427920, 0.5351310, 0.2744800, 0.6231850, 0.8082390, 0.0145753, 0.0308151, 0.7098260, 0.3351360, 0.0502053, 0.3454800, 0.5312370, 0.6644870, 0.8427000, 0.1362940, 0.8458380, 0.0985646, 0.4413880, 0.0276075, 0.6922990, 0.2732090, 0.2214250, 0.0484464, 0.8313440, 0.3083820, 0.6637230, 0.0136811, 0.1782870, 0.2237140, 0.8600840, 0.6575980, 0.9622680, 0.0206604, 0.9074050, 0.7519870, 0.1429680, 0.8462820, 0.1149900, 0.5861740, 0.3372270, 0.2380660, 0.9029480, 0.1271260, 0.7567420, 0.0473744, 0.6056310, 0.3804220, 0.6762140, 0.7460430, 0.5533700, 0.8932570, 0.6069350, 0.1867890, 0.1929530, 0.9506930, 0.9955470, 0.0981962, 0.3909630, 0.7807010, 0.5191070, 0.4965860, 0.7663490, 0.1553120, 0.3047020, 0.2241180, 0.3132420, 0.0265443, 0.9199640, 0.1716210, 0.2551130, 0.1232970, 0.4403120, 0.9618080, 0.4118850, 0.7653890, 0.4068260, 0.7397540, 0.9176630, 0.5442630, 0.1735290, 0.4178260, 0.6174230, 0.8238140, 0.0160507, 0.4372960, 0.7267680, 0.8464350, 0.9754660, 0.3021700, 0.2642090, 0.4599860, 0.3356850, 0.2272060, 0.7274470, 0.6600660, 0.1121980, 0.2116870, 0.6525280, 0.0090506, 0.7118230, 0.1943640, 0.3319040, 0.0903404, 0.8770610, 0.0296722, 0.6993970, 0.8926280, 0.6003860, 0.4938620, 0.4721590, 0.0939505, 0.9182450, 0.1843060, 0.0163192, 0.3436810, 0.2618140, 0.6480670, 0.6516530, 0.2695460, 0.9261880, 0.4803880, 0.4344930, 0.3993830, 0.2461050, 0.5923940, 0.8630590, 0.7871650, 0.0476970, 0.5295820, 0.5576860, 0.2022010, 0.8708390, 0.6478910, 0.7113620, 0.9857960, 0.3253280, 0.7202120, 0.4622890, 0.2539320, 0.4390250, 0.6964840, 0.5769760, 0.4853910, 0.6607030, 0.7361360, 0.1992350, 0.8118550, 0.1123720, 0.8881700, 0.2353430, 0.2113720, 0.1234910, 0.1383800, 0.4780940, 0.3551650, 0.0553904, 0.4594260, 0.3652790, 0.3981480, 0.6998920, 0.5335210, 0.9273590, 0.7369100, 0.8075120, 0.4069940, 0.3834170, 0.1224760, 0.4230170, 0.4634270, 0.6544820, 0.6627390, 0.5836110, 0.1651200, 0.1123640, 0.8766970, 0.5895210, 0.5473410, 0.2438730, 0.9441410, 0.4942600, 0.6139310, 0.8839550, 0.7232270, 0.6323600, 0.3966890, 0.2703390, 0.8261850, 0.0528625, 0.9462030, 0.8448450, 0.3210000, 0.2904950, 0.4259050, 0.6869460, 0.2426460, 0.3800390, 0.7048710, 0.3032290, 0.3572190, 0.3185930, 0.9593820, 0.9233860, 0.8214750, 0.3135930, 0.7171920, 0.4810410, 0.4639540, 0.1152750, 0.3513680, 0.0853185, 0.7940250, 0.5885360, 0.5443030, 0.8920630, 0.3640370, 0.6712570, 0.5936040, 0.5974110, 0.1523290, 0.1288330, 0.4057160, 0.6412140, 0.7097490, 0.7724180, 0.1461600, 0.3118090, 0.5021830, 0.9583850, 0.4886900, 0.0857153, 0.4132520, 0.1028070, 0.9610070, 0.1481840, 0.2482880, 0.7996820, 0.0772276, 0.3534530, 0.0887635, 0.9500900, 0.6728050, 0.4108150, 0.3044310, 0.0617629, 0.5760760, 0.2418140, 0.7278980, 0.5694120, 0.7416550, 0.8676110, 0.5256520, 0.5616740, 0.6006330, 0.1513160, 0.5849320, 0.1662010, 0.4797030, 0.7578830, 0.8930110, 0.3152040, 0.7798220, 0.8953640, 0.7958820, 0.7857110, 0.4659250, 0.8734200, 0.1246710, 0.1992820, 0.7214200, 0.4007280, 0.9972330, 0.7213550, 0.1124510, 0.1080360, 0.7633730, 0.7162330, 0.3347800, 0.9269300, 0.0225535, 0.8067450, 0.0297572, 0.9192840, 0.5893520, 0.3610420, 0.0493033, 0.7463380, 0.1623840, 0.4748220, 0.9601690, 0.1172190, 0.5450770, 0.3230050, 0.5636880, 0.7945650, 0.0392132, 0.6880240, 0.6290370, 0.6506470, 0.3054840, 0.6620050, 0.3484310, 0.8552850, 0.6720880, 0.3311170, 0.2407680, 0.0865616, 0.0736652, 0.3783230, 0.9028160, 0.8407010, 0.9054940, 0.8772190, 0.8519280, 0.0393292, 0.0658117, 0.4320370, 0.0589811, 0.4380080, 0.1634660, 0.2810260, 0.4393540, 0.3617530, 0.5196020, 0.2074950, 0.9293180, 0.8025690, 0.2352560, 0.4827380, 0.1577560, 0.2662830, 0.5181630, 0.0021028, 0.6448530, 0.5546660, 0.0119231, 0.8193530, 0.6457250, 0.3117510, 0.2461400, 0.1773260, 0.2948360, 0.5303500, 0.2642080, 0.0724153, 0.4652490, 0.2932670, 0.4105000, 0.6537910, 0.3520320, 0.8043360, 0.0108138, 0.2585310, 0.8788760, 0.6408150, 0.2785780, 0.9532210, 0.3862290, 0.2672570, 0.8311480, 0.7055500, 0.5460020, 0.5357850, 0.4225280, 0.6789940, 0.7252410, 0.7949890, 0.8520590, 0.8166540, 0.5447130, 0.5587090, 0.1954530, 0.3529600, 0.6858700, 0.2556020, 0.6755060, 0.2288860, 0.4486360, 0.0272089, 0.0022587, 0.3816500, 0.9903850, 0.5606050, 0.7847000, 0.3474850, 0.5552120, 0.7528180, 0.6799050, 0.6893500, 0.4675850, 0.1762070, 0.1158220, 0.5679270, 0.2094570, 0.5527700, 0.4260130, 0.7752620, 0.1750350, 0.5730380, 0.6168700, 0.8256110, 0.7715150, 0.5675050, 0.9558340, 0.3398100, 0.4179650, 0.5188010, 0.6122670, 0.1746520, 0.8565830, 0.6240660, 0.6124420, 0.2110160, 0.9583780, 0.8427820, 0.7312430, 0.1655330, 0.8021940, 0.4256610, 0.4095320, 0.7539400, 0.5273180, 0.2380530, 0.6320160, 0.6499570, 0.5562390, 0.6576140, 0.9749390, 0.1020130, 0.0716261, 0.0773004, 0.8643320, 0.9330250, 0.5314740, 0.1908880, 0.1213480, 0.5011900, 0.0668750, 0.4210410, 0.7096520, 0.1063460, 0.7797000, 0.8489460, 0.1157420, 0.2920940, 0.0250468, 0.5508310, 0.3168480, 0.5226650, 0.9017160, 0.1136490, 0.5944650, 0.8194280, 0.3682170, 0.5607370, 0.3083550, 0.7484350, 0.1539070, 0.5460180, 0.9788920, 0.5673470, 0.9535720, 0.5390740, 0.0806195, 0.8049990, 0.4655740, 0.0566749, 0.6961340, 0.8163100, 0.2667250, 0.5222690, 0.1017640, 0.1789460, 0.1283940, 0.2850240, 0.4091790, 0.6348500, 0.8344920, 0.8145970, 0.5105730, 0.7199740, 0.6053420, 0.0341482, 0.7731870, 0.7246160, 0.5783060, 0.0421734, 0.4355150, 0.9788750, 0.0227986, 0.3063410, 0.2946120, 0.1944230, 0.8080350, 0.9663310, 0.7071180, 0.9129450, 0.4167470, 0.3288750, 0.8756650, 0.6072190, 0.6386120, 0.3054070, 0.0875608, 0.3169390, 0.9278210, 0.1948870, 0.9783080, 0.2685920, 0.7883400, 0.6633210, 0.9630090, 0.6424230, 0.0514480, 0.0534941, 0.7212670, 0.2372750, 0.8847450, 0.7359590, 0.4180720, 0.9576880, 0.5645850, 0.2531380, 0.9454010, 0.3023940, 0.7352810, 0.3074710, 0.2598790, 0.1957900, 0.5137790, 0.0648751, 0.6415900, 0.2309340, 0.6125980, 0.7612530, 0.4798190, 0.4873390, 0.4615880, 0.9078320, 0.1083870, 0.9553460, 0.1361340, 0.1596670, 0.6685840, 0.1409410, 0.9396640, 0.4348990, 0.0029462, 0.6658180, 0.9366360, 0.3175990, 0.9606250, 0.5333840, 0.4780970, 0.7832810, 0.6361920, 0.0692680, 0.1013650, 0.5440360, 0.5515610, 0.4353770, 0.8567990, 0.8644370, 0.8087910, 0.8433500, 0.5823780, 0.1161190, 0.3237340, 0.5794230, 0.6810030, 0.4165300, 0.9785400, 0.9871170, 0.9920680, 0.0712266, 0.8832600, 0.5324630, 0.3068490, 0.1965110, 0.7742080, 0.2624970, 0.3334800, 0.4520720, 0.2436870, 0.7241510, 0.2534170, 0.3279670, 0.3142070, 0.8281360, 0.6684530, 0.8092360, 0.4405780, 0.8006890, 0.1463710, 0.9376490, 0.7661530, 0.0799064, 0.9833990, 0.8828940, 0.3066710, 0.0636027, 0.7356330, 0.3319320, 0.6955190, 0.3403970, 0.2001120, 0.5667220, 0.0527279, 0.7467180, 0.6673630, 0.6241570, 0.6190990, 0.7338490, 0.1438910, 0.5941860, 0.1616130, 0.8647420, 0.6813030, 0.6907640, 0.4774860, 0.2018890, 0.2527850, 0.2816470, 0.7274120, 0.4349930, 0.0033240, 0.9840230, 0.6985930, 0.3936870, 0.6034820, 0.0267820, 0.1800390, 0.9567710, 0.8111580, 0.5176030, 0.0020795, 0.2076320, 0.4471120, 0.2244650, 0.3171290, 0.5184360, 0.7068580, 0.7424410, 0.8601540, 0.7454270, 0.3347630, 0.2691640, 0.4944490, 0.8378000, 0.1272540, 0.3015230, 0.2228080, 0.2824750, 0.5625070, 0.1227960, 0.1154260, 0.5441830, 0.2814370, 0.8023340, 0.7260970, 0.0534124, 0.8909270, 0.3491170, 0.6924500, 0.0812723, 0.0793325, 0.9732190, 0.9797520, 0.3101220, 0.3760030, 0.6669030, 0.0817827, 0.5238490, 0.8284050, 0.8627320, 0.4513120, 0.8214450, 0.4121840, 0.1185350, 0.8058710, 0.4077760, 0.8800920, 0.5693660, 0.8244080, 0.6279010, 0.3477610, 0.0170515, 0.9204380, 0.0083317, 0.0366387, 0.4498070, 0.1936300, 0.5425140, 0.5485160, 0.8161980, 0.4474990, 0.7766600, 0.9853360, 0.6561740, 0.1033500, 0.7550380, 0.1774850, 0.5613510, 0.8613720, 0.2300320, 0.3345730, 0.8077460, 0.3733480, 0.5896040, 0.6708990, 0.0481772, 0.2793580, 0.3050500, 0.5256890, 0.4093550, 0.0005477, 0.7885260, 0.2480070, 0.1068680, 0.4001310, 0.7258190, 0.9810370, 0.4391610, 0.5322690, 0.9896010, 0.2572800, 0.4492730, 0.2475980, 0.7802730, 0.7702510, 0.6366280, 0.6412730, 0.4232470, 0.9565140, 0.9114910, 0.3959000, 0.0769485, 0.0454260, 0.7219510, 0.8643700, 0.6896850, 0.2601620, 0.9074520, 0.1220960, 0.3287040, 0.4965680, 0.1369210, 0.8438760, 0.8011020, 0.3607010, 0.5630070, 0.6268900, 0.2831540, 0.2173900, 0.7253110, 0.8551660, 0.5586560, 0.9673580, 0.9643780, 0.4494300, 0.8731710, 0.3017610, 0.6494250, 0.6467280, 0.2290320, 0.6016050, 0.4087090, 0.7658220, 0.3952470, 0.9751870, 0.8726220, 0.1306720, 0.4461120, 0.1758550, 0.3265190, 0.3809800, 0.0309117, 0.1779660, 0.9905510, 0.9078800, 0.8748140, 0.7844230, 0.1815610, 0.5073550, 0.2375980, 0.6130850, 0.6163960, 0.6309500, 0.1593420, 0.4773830, 0.6187250, 0.4403240, 0.9566730, 0.8861390, 0.6206860, 0.7980950, 0.1188330, 0.0366834, 0.0517451, 0.1437300, 0.4301520, 0.1998630, 0.8170750, 0.5704160, 0.7727970, 0.8625350, 0.6605640, 0.1911100, 0.0655730, 0.6913140, 0.7175620, 0.7422450, 0.5409670, 0.6483250, 0.8100160, 0.2299750, 0.6237020, 0.7076150, 0.3377250, 0.7237570, 0.7484150, 0.8937430, 0.1858000, 0.0539425, 0.0153412, 0.5450980, 0.6192850, 0.1765900, 0.5435690, 0.3955420, 0.5707050, 0.2540370, 0.8722210, 0.6007570, 0.9787890, 0.8038730, 0.2017860, 0.5024590, 0.9305580, 0.7334050, 0.3162430, 0.2057090, 0.9583060, 0.0455077, 0.5739440, 0.3403770, 0.4697360, 0.8854090, 0.8613010, 0.6121920, 0.8769720, 0.3117500, 0.5473290, 0.6468770, 0.7259630, 0.0521066, 0.3740770, 0.9770100, 0.5180610, 0.7506420, 0.5720420, 0.6643400, 0.6901240, 0.2271520, 0.6275120, 0.8265370, 0.9065470, 0.3792270, 0.4321430, 0.2772860, 0.4633460, 0.6364670, 0.9755050, 0.2770730, 0.3676710, 0.5592750, 0.7172140, 0.3604880, 0.6094600, 0.3359190, 0.3537050, 0.6564570, 0.2804880, 0.7670370, 0.3615240, 0.5298610, 0.1318140, 0.6547340, 0.7347130, 0.5875180, 0.8675100, 0.5547600, 0.9693780, 0.5786810, 0.4573410, 0.7800020, 0.3351970, 0.8276630, 0.1343980, 0.0630840, 0.7606170, 0.0676292, 0.6738250, 0.8484020, 0.7197910, 0.1803000, 0.2321630, 0.6237690, 0.4833650, 0.5170620, 0.6174090, 0.8671570, 0.5104470, 0.5638360, 0.0539236, 0.9926290, 0.1892250, 0.3809680, 0.6361420, 0.5574330, 0.3156440, 0.5216740, 0.1756760, 0.4359630, 0.0085285, 0.1473080, 0.7936600, 0.1693800, 0.3459480, 0.2115620, 0.5121720, 0.6811030, 0.6972290, 0.4036110, 0.2912160, 0.4488170, 0.8782500, 0.2642840, 0.7338440, 0.3293910, 0.2199590, 0.0260101, 0.0648996, 0.9086000, 0.0346680, 0.5646310, 0.5142060, 0.7214460, 0.7500700, 0.2172890, 0.7672070, 0.8112160, 0.3703990, 0.0196535, 0.0446292, 0.9948220, 0.0247361, 0.8773000, 0.3872070, 0.0820872, 0.6101540, 0.8883640, 0.0462675, 0.1079090, 0.5165780, 0.0088942, 0.4602930, 0.0035386, 0.2053120, 0.3703430, 0.8264160, 0.8279990, 0.7114610, 0.3888120, 0.2536870, 0.7473450, 0.5543370, 0.2069670, 0.9858840, 0.6273680, 0.9011900, 0.4628030, 0.5189500, 0.4094520, 0.7573360, 0.9804400, 0.9515850, 0.2716240, 0.4601510, 0.2282840, 0.1427380, 0.9249820, 0.4170030, 0.4269810, 0.5601620, 0.1116410, 0.1494830, 0.8947900, 0.7539810, 0.2778950, 0.4576020, 0.0544319, 0.8316430, 0.2834310, 0.8441070, 0.2740680, 0.4665980, 0.5546800, 0.2202460, 0.8596360, 0.1823280, 0.8924850, 0.8778510, 0.6988560, 0.8027100, 0.6197840, 0.5581090, 0.3781950, 0.1266920, 0.4674370, 0.7961670, 0.2383050, 0.6803540, 0.9545010, 0.1337580, 0.3140320, 0.5799850, 0.3041770, 0.9466510, 0.9740110, 0.5264010, 0.7854080, 0.9781460, 0.1471390, 0.4101480, 0.0532675, 0.5461940, 0.7846910, 0.5068830, 0.5323410, 0.4553830, 0.9786530, 0.6051610, 0.0687639, 0.6960010, 0.1796680, 0.2604050, 0.0542478, 0.1299710, 0.1262760, 0.2196100, 0.9177930, 0.6636220, 0.2048640, 0.4838380, 0.9990000, 0.6594930, 0.8021310, 0.6706780, 0.2280720, 0.1903070, 0.9392380, 0.9562390, 0.1795930, 0.4880790, 0.0571219, 0.8481920, 0.3315420, 0.3989840, 0.5815100, 0.8963800, 0.4294670, 0.6120300, 0.4393930, 0.0531025, 0.4424720, 0.8848820, 0.3405080, 0.6216000, 0.5324030, 0.8351120, 0.0589898, 0.6366580, 0.5296830, 0.3443790, 0.8746830, 0.2953320, 0.6777860, 0.6128520, 0.5737530, 0.3345750, 0.8262290, 0.2237820, 0.0354772, 0.4643070, 0.1151680, 0.2120820, 0.9820590, 0.7684740, 0.9393170, 0.9187690, 0.7003480, 0.0988068, 0.5768130, 0.6642750, 0.2193730, 0.0295782, 0.8539600, 0.6450140, 0.0708337, 0.8583090, 0.8069470, 0.0177462, 0.8564830, 0.1572390, 0.4393830, 0.4779610, 0.9927320, 0.9994940, 0.1325290, 0.5126700, 0.0286984, 0.4418010, 0.9749670, 0.9909170, 0.4823330, 0.1005270, 0.0246981, 0.6540180, 0.5183490, 0.1666760, 0.4466020, 0.8712280, 0.1572160, 0.1116460, 0.2290370, 0.0872915, 0.0376411, 0.1127990, 0.6759860, 0.4896300, 0.2178320, 0.2233350, 0.1935630, 0.7982440, 0.8013010, 0.5112020, 0.1294090, 0.8417580, 0.4232530, 0.1284690, 0.7321450, 0.7805980, 0.6908720, 0.1046180, 0.0371630, 0.2470540, 0.0478596, 0.7194050, 0.8704840, 0.3542580, 0.7580100, 0.2531110, 0.4025140, 0.8736540, 0.5634170, 0.9993780, 0.0304160, 0.3413000, 0.7622720, 0.7221460, 0.9047910, 0.1684630, 0.7385260, 0.0282286, 0.4818130, 0.1923580, 0.2268580, 0.9907020, 0.5279990, 0.1194200, 0.0193656, 0.3973230, 0.5924390, 0.1985990, 0.6721430, 0.1752360, 0.3908170, 0.1170820, 0.5604350, 0.0580966, 0.2644960, 0.2834320, 0.7657920, 0.4667030, 0.2020860, 0.4516720, 0.3433530, 0.7264820, 0.4415310, 0.9118900, 0.0299803, 0.3933070, 0.3876230, 0.8299340, 0.3075650, 0.4818080, 0.6667820, 0.1749140, 0.8246550, 0.1378240, 0.9315710, 0.7094690, 0.9728320, 0.4451540, 0.3242200, 0.9008540, 0.9936550, 0.3954040, 0.5710750, 0.5166470, 0.1214790, 0.7505520, 0.8829130, 0.1447570, 0.9862320, 0.6961890, 0.7692760, 0.6249810, 0.4692120, 0.8236870, 0.4897880, 0.7852480, 0.2837160, 0.3229370, 0.7362330, 0.6478940, 0.2877760, 0.5491580, 0.1646500, 0.4893980, 0.2251970, 0.1935530, 0.3360000, 0.0469130, 0.7932840, 0.9790750, 0.3304650, 0.2747080, 0.8129940, 0.5991150, 0.8061250, 0.7380590, 0.2175490, 0.5347880, 0.1575990, 0.1059060, 0.5825820, 0.2667360, 0.3425130, 0.3706090, 0.9618980, 0.8153730, 0.5945240, 0.4376960, 0.4470950, 0.7024700, 0.6023110, 0.5908010, 0.4947400, 0.3739790, 0.5793250, 0.1010750, 0.0626308, 0.3370290, 0.6698180, 0.1628280, 0.8733500, 0.9173020, 0.5056530, 0.8362480, 0.1920470, 0.1952730, 0.5886010, 0.8590410, 0.6530210, 0.6924380, 0.5607650, 0.4077230, 0.0888104, 0.2161150, 0.4566780, 0.1612800, 0.0260849, 0.2998790, 0.8882270, 0.7271020, 0.8702040, 0.4298710, 0.7151670, 0.3084200, 0.6896100, 0.4916560, 0.8386460, 0.7487190, 0.6400050, 0.3979110, 0.0897753, 0.5684690, 0.5126530, 0.9833560, 0.7786310, 0.1051840, 0.6592440, 0.9823780, 0.4743110, 0.4596700, 0.4121080, 0.3900170, 0.8837010, 0.6400170, 0.9320580, 0.7899870, 0.1426160, 0.3365590, 0.8205950, 0.3144310, 0.1269360, 0.4399530, 0.2408670, 0.3123640, 0.7188090, 0.4120390, 0.8171820, 0.3219030, 0.4496370, 0.4035080, 0.1493370, 0.4090090, 0.0146631, 0.6618680, 0.3275440, 0.3159390, 0.2181340, 0.0966501, 0.5730500, 0.5481860, 0.9990180, 0.1550770, 0.6633870, 0.8919640, 0.2811230, 0.9788560, 0.3442500, 0.3306210, 0.9996170, 0.7505080, 0.7052190, 0.6901530, 0.9564010, 0.4998820, 0.8624010, 0.7010780, 0.3994700, 0.9951170, 0.7322610, 0.3183580, 0.9059580, 0.0563059, 0.4960120, 0.2489680, 0.9512360, 0.9704380, 0.4259370, 0.3846900, 0.5031830, 0.2241310, 0.2355360, 0.2324630, 0.1134820, 0.3146160, 0.5832480, 0.5452200, 0.0050315, 0.3363320, 0.1590830, 0.7887920, 0.4671330, 0.9730500, 0.1720540, 0.3635830, 0.6242940, 0.7816990, 0.6052560, 0.9816140, 0.6485600, 0.0871668, 0.0351374, 0.2634610, 0.8038450, 0.5053380, 0.2588770, 0.0474700, 0.7892790, 0.0645482, 0.8492800, 0.4724500, 0.8377640, 0.7753680, 0.5362410, 0.3254560, 0.5505520, 0.1031760, 0.3952390, 0.9041930, 0.5460460, 0.4273300, 0.6170550, 0.9971660, 0.5819850, 0.4877060, 0.8662220, 0.8810280, 0.4845290, 0.3827190, 0.3529510, 0.5681150, 0.6234830, 0.1034020, 0.9646330, 0.9988480, 0.1632340, 0.8300190, 0.8600730, 0.6399730, 0.6758720, 0.7381690, 0.3971240, 0.0115889, 0.0735703, 0.2860470, 0.7512240, 0.0949597, 0.4779880, 0.3567860, 0.1013950, 0.2162030, 0.1329060, 0.2560560, 0.5020550, 0.2548790, 0.6697490, 0.0957924, 0.8096220, 0.2327970, 0.5626370, 0.7450410, 0.7622650, 0.2886320, 0.0265395, 0.7787620, 0.8672360, 0.0003430, 0.9933210, 0.4910110, 0.7781580, 0.2419400, 0.7902620, 0.8648110, 0.4858940, 0.7610470, 0.7553380, 0.2938790, 0.6711810, 0.4897920, 0.3284010, 0.7634600, 0.7785890, 0.6421220, 0.7085170, 0.6451830, 0.0233633, 0.6131190, 0.8592650, 0.3609450, 0.2660100, 0.8757570, 0.9059190, 0.6542220, 0.3979750, 0.1952720, 0.1897350, 0.7892550, 0.7830830, 0.0527582, 0.8749510, 0.4224070, 0.7612440, 0.1699140, 0.5708830, 0.8094120, 0.8563170, 0.8350500, 0.5667220, 0.6154470, 0.9454090, 0.6257340, 0.9397030, 0.4090020, 0.8321190, 0.5678710, 0.3872360, 0.3981200, 0.7531100, 0.5586960, 0.3350570, 0.9322540, 0.5378600, 0.3800240, 0.6142740, 0.7957460, 0.8715340, 0.5132730, 0.1011020, 0.6960520, 0.4055020, 0.2892720, 0.6206970, 0.3973380, 0.5058480, 0.8377330, 0.5107750, 0.6119940, 0.4287680, 0.1297980, 0.7651990, 0.4342630, 0.7731070, 0.5224750, 0.7536500, 0.8040260, 0.9317690, 0.8329120, 0.0880504, 0.2056390, 0.4115860, 0.1083340, 0.4264850, 0.0411395, 0.3607130, 0.8254800, 0.0989515, 0.8331560, 0.3605000, 0.5215620, 0.5281310, 0.8636070, 0.1934740, 0.1629780, 0.2193060, 0.7270790, 0.2783090, 0.0869119, 0.6487460, 0.0426521, 0.0000356, 0.5290620, 0.6048800, 0.8574590, 0.8780030, 0.6053870, 0.4019650, 0.4670080, 0.6107720, 0.0709958, 0.1454140, 0.4443560, 0.9948260, 0.6884880, 0.6762430, 0.9605530, 0.8024740, 0.3255920, 0.1930690, 0.4787500, 0.7101060, 0.9214300, 0.7841020, 0.7801280, 0.1000340, 0.3966610, 0.6353700, 0.5045450, 0.5500060, 0.3479270, 0.6389160, 0.8152630, 0.7294890, 0.1002510, 0.6124880, 0.4600540, 0.8674830, 0.2391040, 0.6000910, 0.6337950, 0.6622010, 0.6117310, 0.2095540, 0.7912280, 0.3605750, 0.6408360, 0.6987910, 0.9366700, 0.5235050, 0.0045225, 0.2973640, 0.6295580, 0.2260650, 0.7317780, 0.0839467, 0.1017700, 0.0606118, 0.9401410, 0.3061260, 0.3451620, 0.5431920, 0.3157550, 0.9511320, 0.4523290, 0.0980958, 0.2802700, 0.8352820, 0.4133150, 0.8847360, 0.0619267, 0.9848360, 0.0044503, 0.1779150, 0.0635478, 0.5682200, 0.3319270, 0.2958940, 0.4100440, 0.5882420, 0.2182290, 0.5846390, 0.6698760, 0.1569730, 0.4918900, 0.8016910, 0.1415090, 0.0675855, 0.0781144, 0.8296450, 0.9140520, 0.9680990, 0.2711510, 0.4060920, 0.7422890, 0.9221060, 0.8663150, 0.1342160, 0.8899120, 0.0267774, 0.7422780, 0.5368520, 0.3102210, 0.4209360, 0.5064550, 0.3929280, 0.3587570, 0.3333610, 0.0968281, 0.4167570, 0.1316190, 0.1931320, 0.1464030, 0.8977020, 0.9628820, 0.8310710, 0.0066635, 0.7360120, 0.0818158, 0.8923810, 0.7065310, 0.2313930, 0.1971580, 0.9305890, 0.6621380, 0.9883440, 0.7690350, 0.4046370, 0.0750083, 0.9517930, 0.7671170, 0.4505650, 0.6518690, 0.7251460, 0.5289000, 0.5318780, 0.4168310, 0.8876740, 0.4088590, 0.9007470, 0.6084170, 0.8959290, 0.7356880, 0.2819830, 0.9907310, 0.4724210, 0.2576640, 0.0528040, 0.9584730, 0.1660910, 0.5380820, 0.7831570, 0.1042970, 0.4260320, 0.4204610, 0.8750190, 0.9985840, 0.9018110, 0.7237670, 0.0864954, 0.7423330, 0.2017040, 0.1858140, 0.3678340, 0.5633030, 0.0655784, 0.6149500, 0.5849770, 0.1786140, 0.0672599, 0.2577030, 0.8445620, 0.9364700, 0.2618600, 0.3742330, 0.8812250, 0.8537060, 0.0870162, 0.3855670, 0.4835590, 0.0128096, 0.4370690, 0.0414377, 0.5790660, 0.7203260, 0.0132674, 0.7203720, 0.1949000, 0.2908990, 0.2982670, 0.8728290, 0.9859840, 0.8563740, 0.3599230, 0.3102500, 0.0663682, 0.6923380, 0.2610270, 0.1095800, 0.0434432, 0.5592150, 0.4140870, 0.9889710, 0.9812720, 0.7227320, 0.3706570, 0.0508580, 0.0109349, 0.3841010, 0.6832770, 0.9433750, 0.7822450, 0.3885320, 0.0053649, 0.4595500, 0.4633200, 0.0019431, 0.8329560, 0.3758310, 0.3341990, 0.2830530, 0.6008680, 0.8801170, 0.8535420, 0.0023379, 0.5855020, 0.9777100, 0.1222090, 0.9653340, 0.6189720, 0.6517940, 0.8601170, 0.4550240, 0.8099910, 0.8122060, 0.6913400, 0.7276350, 0.3167670, 0.5314190, 0.4382140, 0.9919010, 0.9418240, 0.7535560, 0.5857600, 0.6566940, 0.8154600, 0.4084360, 0.7296190, 0.8749690, 0.2296700, 0.7061340, 0.6086140, 0.2700960, 0.8304370, 0.3746840, 0.8633800, 0.0969187, 0.6651930, 0.0514765, 0.7890340, 0.2464760, 0.6864850, 0.9024960, 0.3316140, 0.8761170, 0.9001950, 0.7718790, 0.5633960, 0.3502450, 0.2673340, 0.7055430, 0.6291240, 0.8071090, 0.5907620, 0.6543370, 0.2574850, 0.1389600, 0.2723420, 0.6430330, 0.6687210, 0.0639907, 0.0826861, 0.1262190, 0.5073710, 0.1703060, 0.1497790, 0.8902350, 0.9334650, 0.2987020, 0.0844281, 0.4729510, 0.7836540, 0.6667880, 0.2024390, 0.9183370, 0.3282400, 0.2166790, 0.7239950, 0.8142900, 0.3431510, 0.4523430, 0.4336870, 0.7438880, 0.9096790, 0.1978770, 0.5076020, 0.5082820, 0.2388350, 0.1944740, 0.1596480, 0.2717620, 0.5302760, 0.5963540, 0.3039220, 0.5672440, 0.1109690, 0.5414500, 0.2569620, 0.1588530, 0.6249430, 0.4153930, 0.7321280, 0.5760830, 0.0521967, 0.1605870, 0.9749150, 0.1774170, 0.0848106, 0.4193280, 0.1782720, 0.0925567, 0.9610990, 0.3940140, 0.1579680, 0.5669410, 0.1605910, 0.7236270, 0.2260130, 0.7926460, 0.7595760, 0.0415816, 0.4095700, 0.3248340, 0.9201240, 0.5016910, 0.7706220, 0.4017740, 0.1250070, 0.8606020, 0.1452310, 0.8502310, 0.2043040, 0.1794050, 0.1689800, 0.0354179, 0.7976200, 0.3214980, 0.7447260, 0.0264040, 0.3122670, 0.4911550, 0.0362320, 0.6455040, 0.6872350, 0.1599830, 0.6529860, 0.1803530, 0.3575440, 0.0612027, 0.0009369, 0.6141880, 0.3706270, 0.1351060, 0.8952340, 0.4551970, 0.1953470, 0.9153400, 0.8584860, 0.9539290, 0.9214880, 0.5219010, 0.3530690, 0.9470570, 0.9132550, 0.2242020, 0.6148870, 0.9398020, 0.0929465, 0.3148370, 0.6310560, 0.2283550, 0.5991050, 0.8567990, 0.0120713, 0.8396700, 0.8915920, 0.7484880, 0.2589910, 0.2501330, 0.3120440, 0.3877810, 0.9622160, 0.2972400, 0.0627565, 0.9935920, 0.3211350, 0.2116090, 0.4577670, 0.5526380, 0.4249470, 0.6197980, 0.7487990, 0.5933190, 0.0857750, 0.5194510, 0.7200460, 0.2452800, 0.6803130, 0.8928120, 0.3777540, 0.6774690, 0.8155570, 0.3418570, 0.5688860, 0.2361400, 0.8987110, 0.5853520, 0.7078230, 0.0714605, 0.2066970, 0.9056360, 0.2725520, 0.2618640, 0.2347240, 0.7928690, 0.9473830, 0.4876450, 0.9504430, 0.0804064, 0.7128080, 0.0780785, 0.7734880, 0.8847070, 0.1148330, 0.4581680, 0.1182280, 0.0087679, 0.2714500, 0.9966670, 0.0650028, 0.8721750, 0.7108120, 0.4029430, 0.6215460, 0.3684850, 0.3118320, 0.5684940, 0.8716160, 0.7494180, 0.0886400, 0.9163690, 0.3236740, 0.3245860, 0.3667240, 0.4234530, 0.5434380, 0.8283440, 0.4117870, 0.9543690, 0.8824780, 0.9180500, 0.2338530, 0.1245400, 0.7499460, 0.2514620, 0.5977860, 0.1002380, 0.5571310, 0.1917850, 0.4564440, 0.5653170, 0.7444370, 0.0781992, 0.4380340, 0.5327560, 0.6415720, 0.9290550, 0.7099770, 0.2655590, 0.2142770, 0.5823430, 0.0437601, 0.7270980, 0.5856020, 0.1943580, 0.9970430, 0.1261080, 0.5062850, 0.5840450, 0.7460320, 0.1592350, 0.9304530, 0.5434870, 0.0672393, 0.5352710, 0.8631800, 0.2763430, 0.6319790, 0.2071610, 0.1585850, 0.4433560, 0.4876940, 0.4135800, 0.1882580, 0.3237580, 0.3846190, 0.0117183, 0.8823970, 0.3542970, 0.1073500, 0.5963280, 0.7514750, 0.9412650, 0.1743120, 0.2829840, 0.2440430, 0.7812980, 0.4483420, 0.2302320, 0.3634900, 0.8382520, 0.6476110, 0.4784550, 0.1969970, 0.4703410, 0.0604516, 0.0472010, 0.9251650, 0.8377970, 0.8210420, 0.8148680, 0.6040560, 0.5033980, 0.2191050, 0.3828250, 0.4119990, 0.8309260, 0.7719620, 0.4639800, 0.3872920, 0.5939130, 0.1203910, 0.2341380, 0.4648400, 0.6870560, 0.3386710, 0.5963970, 0.3041090, 0.1601240, 0.7055250, 0.4426190, 0.8356040, 0.9095920, 0.2531330, 0.5644260, 0.5255220, 0.0236053, 0.5980180, 0.1791000, 0.1614100, 0.7484080, 0.5735900, 0.3636730, 0.2475820, 0.2756270, 0.7092460, 0.5890670, 0.5796010, 0.5350830, 0.0376110, 0.7718190, 0.1796160, 0.6044830, 0.5387660, 0.2690970, 0.8041750, 0.2839700, 0.3865580, 0.8134650, 0.1242400, 0.1808260, 0.3350990, 0.8467160, 0.3770300, 0.4685060, 0.5398670, 0.8215430, 0.6518680, 0.1933130, 0.3077620, 0.7901540, 0.2734400, 0.4866450, 0.3915520, 0.5063640, 0.5377500, 0.6319740, 0.8668110, 0.6274370, 0.6568830, 0.9165150, 0.2767810, 0.8768590, 0.8516320, 0.6289110, 0.2762630, 0.7551390, 0.3983020, 0.3172850, 0.9657450, 0.5396790, 0.3864950, 0.8680920, 0.9072110, 0.0888999, 0.3145080, 0.4413720, 0.2589050, 0.1244320, 0.6234190, 0.1804660, 0.8944920, 0.5592180, 0.0646865, 0.4954880, 0.6079130, 0.7250820, 0.2473890, 0.8357780, 0.4003160, 0.1695250, 0.0871621, 0.7824410, 0.0546528, 0.4536140, 0.3106770, 0.6909020, 0.2852090, 0.0630503, 0.6095540, 0.1778640, 0.5876260, 0.3221260, 0.0634543, 0.3906730, 0.0904105, 0.1787900, 0.9229630, 0.2268270, 0.0848163, 0.3557290, 0.2853850, 0.9386150, 0.0774163, 0.1805110, 0.4560020, 0.1082600, 0.2078100, 0.8761730, 0.2022120, 0.1580890, 0.2476930, 0.3143160, 0.0712029, 0.5952490, 0.5236080, 0.9976040, 0.2293930, 0.8111060, 0.5879310, 0.0965318, 0.6948200, 0.1580200, 0.3612670, 0.2949250, 0.1338840, 0.9338450, 0.2916670, 0.8674210, 0.5022520, 0.4506410, 0.8637050, 0.6069620, 0.4591050, 0.3298180, 0.4061970, 0.4685330, 0.7423880, 0.7617960, 0.5337130, 0.7293590, 0.2822000, 0.9392180, 0.8340020, 0.1212110, 0.6544120, 0.0895728, 0.1170870, 0.9721340, 0.4387620, 0.7893890, 0.5158910, 0.3425840, 0.5282650, 0.6691060, 0.5107200, 0.4492410, 0.3136970, 0.4771140, 0.4161730, 0.6616460, 0.1710660, 0.1930530, 0.5268210, 0.3018690, 0.3002050, 0.1903510, 0.2421930, 0.4666460, 0.5948550, 0.0568293, 0.8525410, 0.7198560, 0.6760350, 0.5892780, 0.5553000, 0.4240110, 0.5178210, 0.4542810, 0.8525500, 0.5063520, 0.9705900, 0.7008180, 0.4213320, 0.2612120, 0.0735979, 0.0027166, 0.5605140, 0.6893450, 0.6148410, 0.7635020, 0.5827230, 0.9558110, 0.4796980, 0.0131003, 0.0843812, 0.7966580, 0.5883490, 0.1558680, 0.6577900, 0.9825380, 0.6718650, 0.1050120, 0.2391210, 0.0077177, 0.0866143, 0.6086780, 0.5580950, 0.9831750, 0.0165262, 0.3576750, 0.0002785, 0.7009730, 0.4951330, 0.8427580, 0.9202550, 0.0947307, 0.6140430, 0.8982900, 0.1469040, 0.3476330, 0.4187200, 0.6612270, 0.5211980, 0.5479090, 0.1628080, 0.8973360, 0.2076760, 0.3292920, 0.0743800, 0.6545250, 0.2502010, 0.8533670, 0.8089860, 0.8292560, 0.2364380, 0.5772550, 0.4345380, 0.7534400, 0.1599580, 0.8731130, 0.0207941, 0.6406300, 0.3951710, 0.5121740, 0.4286750, 0.9253810, 0.7996580, 0.3107990, 0.5666870, 0.4028320, 0.0778359, 0.8950300, 0.5827620, 0.6137680, 0.4741980, 0.0009734, 0.2203830, 0.8195020, 0.2264120, 0.3718630, 0.9184790, 0.3537760, 0.1089290, 0.3865100, 0.3189000, 0.7101360, 0.4965680, 0.3145920, 0.5974610, 0.1133250, 0.5465220, 0.1145390, 0.1666220, 0.4142590, 0.1741320, 0.7010650, 0.4105650, 0.4775120, 0.9657650, 0.2404220, 0.4771000, 0.7636310, 0.1366340, 0.1972250, 0.3830500, 0.6893880, 0.9746160, 0.9175830, 0.7911030, 0.7027080, 0.1957880, 0.2793490, 0.1733310, 0.2317190, 0.7373910, 0.1087680, 0.6180880, 0.8572400, 0.6548530, 0.1427330, 0.6815600, 0.2502390, 0.5146000, 0.3372890, 0.0602933, 0.4839390, 0.6873750, 0.9108790, 0.3947470, 0.3822090, 0.8715570, 0.5118430, 0.3883070, 0.6297970, 0.0488000, 0.7562710, 0.9128220, 0.4610640, 0.0126493, 0.8146880, 0.4895760, 0.0651276, 0.5629940, 0.4605340, 0.0348916, 0.6267410, 0.3758820, 0.6677570, 0.1876950, 0.2517230, 0.6108390, 0.3401130, 0.4825160, 0.1303920, 0.8451170, 0.1304770, 0.0247904, 0.8265660, 0.6983100, 0.5068050, 0.0187975, 0.6573940, 0.4771500, 0.2685920, 0.5200650, 0.5330090, 0.4834110, 0.4522240, 0.5730600, 0.1464720, 0.4825910, 0.2169640, 0.3909610, 0.4539200, 0.1175840, 0.9281900, 0.3607660, 0.0496142, 0.5274240, 0.3691490, 0.2952950, 0.4904580, 0.8872960, 0.8159670, 0.8929460, 0.0162312, 0.0848181, 0.0767815, 0.1671990, 0.3596050, 0.1820550, 0.4529730, 0.2884630, 0.6427960, 0.0846377, 0.1173940, 0.5758610, 0.3623400, 0.9717050, 0.7477610, 0.6199640, 0.1468190, 0.3782070, 0.3241240, 0.5760790, 0.7650960, 0.7362280, 0.0579590, 0.0426969, 0.1473200, 0.2903630, 0.3298670, 0.3736300, 0.5389300, 0.7116550, 0.0884120, 0.0707983, 0.2568710, 0.6499040, 0.1405200, 0.3081270, 0.3009490, 0.9756140, 0.6286930, 0.0443345, 0.0250528, 0.4916510, 0.7642410, 0.8506610, 0.6429150, 0.6473070, 0.0055906, 0.5912520, 0.0131474, 0.9010870, 0.2100530, 0.7866630, 0.2648670, 0.9277680, 0.3509240, 0.9524800, 0.8772820, 0.9155740, 0.2437520, 0.9751550, 0.5556150, 0.0290126, 0.3609650, 0.4768730, 0.1175960, 0.8038910, 0.5187840, 0.0200459, 0.8456130, 0.0643111, 0.2712260, 0.1850800, 0.3441180, 0.7036400, 0.2296510, 0.7618570, 0.0952546, 0.1115350, 0.7265590, 0.8670470, 0.8209920, 0.2596790, 0.6180270, 0.1549210, 0.5854770, 0.6060950, 0.9807980, 0.7633490, 0.8045200, 0.8729550, 0.2784620, 0.5050710, 0.9671210, 0.6182230, 0.0693947, 0.6835270, 0.0750411, 0.9239490, 0.2756550, 0.7155360, 0.6369080, 0.5817270, 0.5563330, 0.4288430, 0.1720270, 0.8058320, 0.4393870, 0.7097570, 0.3997130, 0.8278310, 0.8279290, 0.3214910, 0.5917700, 0.4136500, 0.4839520, 0.1903680, 0.0175991, 0.9823740, 0.9184780, 0.8375690, 0.2332290, 0.5499000, 0.7744480, 0.7798170, 0.2559760, 0.5853070, 0.5061700, 0.3034460, 0.9929470, 0.2947630, 0.1562290, 0.3772050, 0.0452779, 0.7364890, 0.4483370, 0.0834545, 0.9790480, 0.9559390, 0.4571810, 0.7871100, 0.4062160, 0.0623600, 0.9564750, 0.3157860, 0.9216230, 0.8219650, 0.8258080, 0.7517210, 0.7758880, 0.7712050, 0.4830520, 0.0400101, 0.0878020, 0.6029270, 0.2799100, 0.8564520, 0.5407250, 0.8127640, 0.1649010, 0.4802610, 0.6442570, 0.9219780, 0.6189890, 0.4376360, 0.5646280, 0.2598990, 0.7550560, 0.0210830, 0.3053250, 0.2197810, 0.7064840, 0.8157460, 0.1466650, 0.2259100, 0.9592090, 0.2996720, 0.9258440, 0.6607470, 0.8804850, 0.3336520, 0.1432840, 0.0752058, 0.4336400, 0.6587820, 0.1474420, 0.9479920, 0.6416510, 0.7837770, 0.4191810, 0.9057130, 0.2173400, 0.7815340, 0.5938680, 0.0403157, 0.2665180, 0.3006280, 0.0222828, 0.2339150, 0.3093490, 0.9322350, 0.1098350, 0.0958970, 0.1702720, 0.2431720, 0.6770870, 0.2350480, 0.1552390, 0.8038240, 0.4419820, 0.0500371, 0.9846520, 0.3397040, 0.8528780, 0.8054580, 0.3825140, 0.2596630, 0.7666920, 0.2303010, 0.8025840, 0.7866460, 0.6980340, 0.8139470, 0.8954000, 0.8588920, 0.8949350, 0.6518520, 0.2407400, 0.0520412, 0.3268660, 0.3688700, 0.8012230, 0.7489080, 0.9217560, 0.4948510, 0.9205770, 0.7356030, 0.9310690, 0.6108890, 0.6190850, 0.7281650, 0.4982990, 0.1566220, 0.2365400, 0.8963310, 0.1755290, 0.8947440, 0.0875276, 0.0224419, 0.3055150, 0.0445080, 0.9910220, 0.4720530, 0.4029860, 0.2781180, 0.2296810, 0.4007420, 0.2694230, 0.5286730, 0.7660470, 0.2104260, 0.7677350, 0.9578210, 0.6247440, 0.5869120, 0.9762290, 0.5752150, 0.5090400, 0.7471480, 0.0752972, 0.1663480, 0.7903760, 0.1207040, 0.7856140, 0.4769160, 0.2118190, 0.8851020, 0.9168510, 0.3465260, 0.3466490, 0.4380510, 0.7776270, 0.7903390, 0.5464350, 0.0126564, 0.5073700, 0.7998920, 0.6355630, 0.5853190, 0.3804820, 0.5174650, 0.0948706, 0.8481480, 0.3338560, 0.1000160, 0.3013890, 0.4141130, 0.0209561, 0.4338820, 0.2443690, 0.1464320, 0.3241480, 0.1411120, 0.9696590, 0.0535825, 0.0686587, 0.7818440, 0.4313660, 0.5643190, 0.1071410, 0.6317520, 0.1433030, 0.6700900, 0.7543650, 0.2912720, 0.1691550, 0.5279260, 0.8343400, 0.2706050, 0.6689800, 0.5794110, 0.4426020, 0.3375140, 0.6858750, 0.1008350, 0.6375170, 0.0208273, 0.1427980, 0.2020160, 0.9112020, 0.1212630, 0.6080150, 0.9301610, 0.4121640, 0.0801841, 0.7425180, 0.6982130, 0.7891510, 0.7421240, 0.6194010, 0.6758710, 0.8138040, 0.8119880, 0.9550540, 0.3139530, 0.1132580, 0.4278080, 0.8070610, 0.7857130, 0.5788650, 0.8365510, 0.5655940, 0.1108930, 0.0327342, 0.5288140, 0.9373530, 0.5954070, 0.4964020, 0.6706470, 0.0111523, 0.6183150, 0.9660890, 0.1617560, 0.3691010, 0.4579260, 0.1873970, 0.5086870, 0.3804510, 0.1013670, 0.3177860, 0.6321020, 0.6399140, 0.7625040, 0.0965030, 0.4433090, 0.4128570, 0.1402940, 0.2731740, 0.8566080, 0.6601650, 0.6576340, 0.4319440, 0.5670710, 0.2604960, 0.9906180, 0.0144212, 0.5940670, 0.2346420, 0.9602980, 0.2097790, 0.9474180, 0.4882820, 0.2458720, 0.2847530, 0.8467170, 0.2999030, 0.2142150, 0.1197060, 0.5965810, 0.7522310, 0.9205600, 0.5881330, 0.9620790, 0.3691430, 0.7436720, 0.3963240, 0.5317920, 0.4403730, 0.9993450, 0.8263950, 0.1538070, 0.6556800, 0.7859500, 0.8094700, 0.0968109, 0.0861839, 0.9994600, 0.1214240, 0.8236140, 0.9102470, 0.8607120, 0.7052450, 0.2423100, 0.3154550, 0.0559218, 0.8596400, 0.4147370, 0.2216810, 0.4736290, 0.8249590, 0.8116890, 0.9375810, 0.4354330, 0.1226930, 0.5265940, 0.5164310, 0.1937840, 0.7320930, 0.1367360, 0.1338750, 0.3816790, 0.8197280, 0.9803640, 0.3644870, 0.9021000, 0.3749950, 0.6041680, 0.9277650, 0.3969680, 0.1101040, 0.5308560, 0.4906450, 0.4627710, 0.7496940, 0.8392610, 0.5644940, 0.8246060, 0.9236210, 0.8483860, 0.1093910, 0.2260180, 0.8070450, 0.4593720, 0.1028680, 0.3586950, 0.8231570, 0.4688060, 0.7281890, 0.6130990, 0.4660010, 0.0035594, 0.2851430, 0.8512640, 0.9737820, 0.8124010, 0.2817710, 0.3619180, 0.6945350, 0.2730440, 0.9303060, 0.1301480, 0.7881210, 0.9575140, 0.1862970, 0.4129950, 0.4409520, 0.0977291, 0.7492240, 0.5920900, 0.5848790, 0.4563070, 0.2329600, 0.2335640, 0.4060920, 0.9413060, 0.0124222, 0.5715120, 0.4351830, 0.1885630, 0.4686630, 0.2180750, 0.4977010, 0.6213190, 0.8724580, 0.7069260, 0.6406800, 0.4305960, 0.0492570, 0.3266790, 0.8301910, 0.2416710, 0.6536480, 0.0506871, 0.8298300, 0.2552790, 0.6383880, 0.7520330, 0.6629430, 0.8260700, 0.7589780, 0.1882630, 0.6585690, 0.4866030, 0.0800300, 0.6441020, 0.3909710, 0.1713940, 0.0401618, 0.1445310, 0.7462190, 0.1662740, 0.3448160, 0.8027020, 0.9575280, 0.0360370, 0.4343550, 0.1426930, 0.5220370, 0.3797390, 0.5980120, 0.6400770, 0.1568110, 0.8902300, 0.6100240, 0.8413840, 0.9917820, 0.0050088, 0.5297500, 0.3008150, 0.9917780, 0.8354790, 0.6498820, 0.6363400, 0.0571184, 0.9119760, 0.1311420, 0.0973227, 0.5645010, 0.3464560, 0.5957290, 0.7019060, 0.7219730, 0.6494840, 0.4175870, 0.1315500, 0.9050520, 0.9825150, 0.8355800, 0.8509280, 0.1535460, 0.5587300, 0.2954100, 0.7658940, 0.1532460, 0.1256430, 0.4444270, 0.0225897, 0.9193360, 0.2992400, 0.6848630, 0.2792180, 0.4025870, 0.8668700, 0.2064260, 0.8230840, 0.1815150, 0.1373330, 0.0429065, 0.2824390, 0.1806980, 0.8223400, 0.8828630, 0.1802530, 0.5356740, 0.8236580, 0.8971740, 0.6506830, 0.8926230, 0.7782570, 0.0859129, 0.1748510, 0.1296230, 0.3616220, 0.0113652, 0.6147430, 0.2735360, 0.1279840, 0.3872540, 0.3198220, 0.3144410, 0.0170322, 0.1918610, 0.4921080, 0.3867410, 0.9500850, 0.7896330, 0.3983300, 0.2002340, 0.1637330, 0.8986660, 0.8543220, 0.1669120, 0.7305190, 0.7032800, 0.2723940, 0.5609200, 0.0120119, 0.9645690, 0.7065630, 0.2512240, 0.1997410, 0.1162890, 0.3509040, 0.5891440, 0.6768390, 0.4192280, 0.8568710, 0.9400850, 0.6619940, 0.4528490, 0.8363960, 0.9669260, 0.5518600, 0.9272070, 0.9749190, 0.4548330, 0.7496490, 0.5729580, 0.3736040, 0.0203335, 0.3947740, 0.4958630, 0.6421280, 0.9696890, 0.5949590, 0.8136900, 0.7378900, 0.5560420, 0.1337570, 0.5502460, 0.8000400, 0.5717710, 0.6604160, 0.4185430, 0.7423490, 0.8033490, 0.2245130, 0.4035770, 0.8442070, 0.0849369, 0.2389580, 0.1289910, 0.0530984, 0.4877150, 0.5394610, 0.5794410, 0.9136440, 0.1599100, 0.3962380, 0.1905950, 0.0924820, 0.4528220, 0.5527650, 0.8166180, 0.4985110, 0.0692012, 0.9805320, 0.3798620, 0.0094907, 0.7161440, 0.8710720, 0.5316720, 0.1360750, 0.7566110, 0.7209060, 0.7188510, 0.9019880, 0.4874330, 0.7723760, 0.1642890, 0.0901189, 0.0412866, 0.8451310, 0.6651940, 0.1924600, 0.7410480, 0.2776750, 0.8814560, 0.0554137, 0.5184730, 0.1521340, 0.3557170, 0.8656810, 0.6345430, 0.4018490, 0.9481040, 0.9010800, 0.5736210, 0.2965430, 0.0763738, 0.7761760, 0.8617760, 0.6372210, 0.5873730, 0.9951020, 0.5112970, 0.6541720, 0.9665040, 0.7211080, 0.6784020, 0.4146450, 0.6843340, 0.9273780, 0.1097660, 0.4731000, 0.5781530, 0.5700030, 0.2514350, 0.7942230, 0.8930170, 0.0516718, 0.0274512, 0.6206690, 0.4592170, 0.6690430, 0.6937990, 0.2370620, 0.8221730, 0.0684886, 0.1854310, 0.3731010, 0.7740470, 0.4719750, 0.4006690, 0.2521690, 0.5398480, 0.2186470, 0.6110290, 0.3159740, 0.3297860, 0.2876630, 0.6415150, 0.4780820, 0.8151850, 0.4868690, 0.3633790, 0.2048510, 0.2380280, 0.0492825, 0.1994460, 0.0204031, 0.2996590, 0.0852887, 0.8946540, 0.2803060, 0.1459910, 0.2853550, 0.9095000, 0.7373800, 0.0975732, 0.2405620, 0.0309165, 0.4566840, 0.8607950, 0.8896140, 0.5771350, 0.2591490, 0.4990090, 0.9005350, 0.7371670, 0.9131560, 0.3655780, 0.5981650, 0.3110320, 0.8416840, 0.0753397, 0.0548202, 0.2236260, 0.1198470, 0.6754960, 0.0390476, 0.2423830, 0.0532638, 0.0861004, 0.4274660, 0.7463400, 0.5827850, 0.1465210, 0.0627763, 0.1581480, 0.5980060, 0.2141650, 0.8806480, 0.3157520, 0.5638260, 0.3270840, 0.5901400, 0.4906820, 0.2706130, 0.5175670, 0.7582430, 0.0910104, 0.7717230, 0.5423790, 0.0631830, 0.4574400, 0.0418066, 0.8203980, 0.5935390, 0.7156740, 0.1340620, 0.0881155, 0.0400552, 0.1171460, 0.9942240, 0.1211620, 0.8191000, 0.3619060, 0.6877200, 0.8144940, 0.3563130, 0.4358670, 0.7108390, 0.5868330, 0.5981820, 0.9806010, 0.6264560, 0.1495580, 0.7077800, 0.9596620, 0.2562770, 0.6966890, 0.3247940, 0.3712300, 0.8616500, 0.3092490, 0.0975485, 0.0131274, 0.9565580, 0.8077770, 0.3538620, 0.0421637, 0.9323790, 0.3106040, 0.0882323, 0.0863957, 0.9118610, 0.5899880, 0.1656960, 0.8151520, 0.4369180, 0.3622640, 0.2401870, 0.8987920, 0.6981300, 0.4174760, 0.0079783, 0.0250784, 0.6655640, 0.9535130, 0.8733050, 0.2833370, 0.5334710, 0.3814030, 0.5673850, 0.1372310, 0.9741000, 0.7818500, 0.3481290, 0.0429646, 0.9205380, 0.2294420, 0.5406940, 0.0548173, 0.8107470, 0.7174830, 0.2380110, 0.5865470, 0.0420907, 0.4848800, 0.8337640, 0.0566183, 0.9579410, 0.3814300, 0.9064690, 0.6194750, 0.6849740, 0.2343470, 0.8199020, 0.9751540, 0.4623000, 0.2361630, 0.3040220, 0.1962120, 0.7811160, 0.0389577, 0.7123150, 0.0646683, 0.3956180, 0.4252860, 0.4312300, 0.7062140, 0.9726520, 0.2862570, 0.3182480, 0.0787501, 0.1204870, 0.6704790, 0.6205500, 0.5670210, 0.9320570, 0.6131380, 0.7091430, 0.8098300, 0.1508120, 0.8311410, 0.6134480, 0.4554930, 0.2504050, 0.5786400, 0.5174960, 0.2309690, 0.2541240, 0.4592140, 0.3099430, 0.0829950, 0.4880020, 0.2392980, 0.9466290, 0.5457690, 0.2239210, 0.9026070, 0.7339960, 0.4961120, 0.7338510, 0.1527010, 0.6368000, 0.9347790, 0.4465630, 0.4084560, 0.6024780, 0.4156750, 0.7489180, 0.9997000, 0.9810320, 0.2790010, 0.6639990, 0.4381390, 0.5805780, 0.6086770, 0.4187310, 0.5188250, 0.6060750, 0.7293540, 0.8603860, 0.0544964, 0.2435410, 0.7616720, 0.7737760, 0.0250009, 0.6265560, 0.9971380, 0.3980050, 0.6453220, 0.3194460, 0.7621710, 0.5220080, 0.5669290, 0.0290330, 0.9726740, 0.7172380, 0.1856570, 0.0426366, 0.3079190, 0.6491140, 0.7968750, 0.9532200, 0.0249678, 0.9126550, 0.8040890, 0.4262210, 0.8098610, 0.3089560, 0.9334720, 0.0102488, 0.1690780, 0.5477650, 0.2805740, 0.3371450, 0.1508840, 0.9357790, 0.1295530, 0.4468520, 0.6659370, 0.4558840, 0.4171390, 0.0346171, 0.0037152, 0.5161320, 0.5609010, 0.8292410, 0.4146880, 0.2425750, 0.8355850, 0.0284572, 0.8349960, 0.1226980, 0.1217590, 0.1205360, 0.1812600, 0.6541520, 0.0024789, 0.8036560, 0.0975604, 0.5312530, 0.2153200, 0.2017920, 0.6427610, 0.9118040, 0.0114661, 0.3147620, 0.3333490, 0.0703683, 0.7502690, 0.5847510, 0.5518250, 0.8201210, 0.9742940, 0.8389790, 0.8313580, 0.3787760, 0.4976070, 0.2601390, 0.9866650, 0.4733350, 0.3006470, 0.4461590, 0.4248710, 0.1771900, 0.2135770, 0.9982520, 0.1747790, 0.9260560, 0.7430900, 0.1813790, 0.0439768, 0.2520420, 0.8043870, 0.2913560, 0.9317090, 0.7465770, 0.9470060, 0.5165500, 0.5854330, 0.0243530, 0.7245040, 0.7684020, 0.4461860, 0.8589190, 0.8823640, 0.0598931, 0.8165510, 0.3831060, 0.0829907, 0.3663920, 0.6749580, 0.5582140, 0.9483420, 0.8638230, 0.2703170, 0.1629110, 0.0368371, 0.3578600, 0.7306200, 0.0788197, 0.5883010, 0.9599290, 0.3690710, 0.3980260, 0.6777220, 0.1885480, 0.8846550, 0.0297477, 0.9352490, 0.8785930, 0.2809460, 0.0187735, 0.5159110, 0.5554580, 0.4119730, 0.3649010, 0.5988810, 0.9872290, 0.3580200, 0.3104880, 0.6927700, 0.3874680, 0.3011050, 0.8350690, 0.3359140, 0.8125800, 0.0380808, 0.0362367, 0.4853040, 0.6508470, 0.3570760, 0.8091500, 0.0491009, 0.4254680, 0.3965070, 0.6634180, 0.1541740, 0.6643210, 0.5568460, 0.7187350, 0.5941260, 0.0746191, 0.1050590, 0.9767730, 0.0889847, 0.0419667, 0.4865160, 0.8833210, 0.4013960, 0.9676930, 0.4816390, 0.9425060, 0.9114930, 0.6405390, 0.5647460, 0.3638980, 0.0607914, 0.5460490, 0.1797110, 0.5819920, 0.0083515, 0.9771950, 0.5285360, 0.6254850, 0.1361570, 0.9305630, 0.1770320, 0.3495030, 0.9479100, 0.5414760, 0.6524910, 0.1634610, 0.7330370, 0.4286700, 0.8567300, 0.7583130, 0.9876680, 0.0093108, 0.4830530, 0.4469710, 0.5245260, 0.5321240, 0.5465640, 0.2917520, 0.5720310, 0.5607350, 0.3288100, 0.0371912, 0.3063460, 0.6189370, 0.8444960, 0.8698090, 0.0505274, 0.0694339, 0.9835740, 0.1110430, 0.6578240, 0.5932200, 0.2613580, 0.2819850, 0.4984390, 0.4112700, 0.3948840, 0.7637640, 0.8138150, 0.8290490, 0.6633190, 0.3230080, 0.7002820, 0.1145920, 0.7162930, 0.4230250, 0.4237710, 0.4355380, 0.7073640, 0.4962320, 0.7264100, 0.6209210, 0.8360250, 0.4693630, 0.5833250, 0.9796160, 0.0983826, 0.5728280, 0.3848140, 0.9255110, 0.0918439, 0.9144780, 0.6478330, 0.1311790, 0.3067650, 0.6677730, 0.4663730, 0.9487780, 0.0436849, 0.5141190, 0.4431280, 0.9952100, 0.6294680, 0.4498490, 0.6675360, 0.2580650, 0.7710280, 0.4164780, 0.8949730, 0.7712660, 0.9344360, 0.0865983, 0.0235080, 0.8898110, 0.1332630, 0.9863740, 0.6155210, 0.0046848, 0.9679490, 0.4220450, 0.2292060, 0.1205970, 0.4434650, 0.9647860, 0.6456510, 0.8792260, 0.1772340, 0.8561580, 0.1398150, 0.7558410, 0.8349670, 0.6979010, 0.1687190, 0.2218660, 0.0547010, 0.6517310, 0.8951550, 0.7953800, 0.9116360, 0.8831500, 0.6975340, 0.6099220, 0.6271220, 0.9615100, 0.3397410, 0.1073180, 0.7892580, 0.6588960, 0.9858180, 0.4897430, 0.8549600, 0.6033880, 0.6926390, 0.3811680, 0.2664050, 0.2541550, 0.3455460, 0.5861160, 0.4457230, 0.3305320, 0.2112650, 0.0306554, 0.7039490, 0.9194060, 0.3640630, 0.1267000, 0.0231864, 0.1543650, 0.9497140, 0.7381610, 0.9679770, 0.3157210, 0.2931990, 0.6816100, 0.5004120, 0.2179230, 0.8668570, 0.7517070, 0.0515239, 0.1500180, 0.6936660, 0.6644300, 0.7354080, 0.4797490, 0.1250810, 0.6552090, 0.2397900, 0.3331880, 0.1327750, 0.8695560, 0.1166860, 0.3747820, 0.1144450, 0.4684000, 0.2682320, 0.9277560, 0.4022780, 0.9644990, 0.5301750, 0.8705400, 0.9655580, 0.0447532, 0.2064610, 0.8107900, 0.3365300, 0.4742400, 0.1910520, 0.3254860, 0.3618800, 0.7198330, 0.3297260, 0.4342730, 0.3230680, 0.8857770, 0.8290580, 0.6118970, 0.1862410, 0.6339040, 0.7685940, 0.1327180, 0.1239320, 0.6359310, 0.9920500, 0.2496100, 0.9404680, 0.1333990, 0.1404370, 0.8590680, 0.6082350, 0.9768010, 0.2029410, 0.7369280, 0.2833890, 0.7142720, 0.5873350, 0.3904340, 0.9859490, 0.9270600, 0.5542910, 0.8345850, 0.7673530, 0.8469630, 0.0895051, 0.5380470, 0.6392030, 0.9246170, 0.9972880, 0.5821030, 0.6891800, 0.4239010, 0.1556800, 0.8903140, 0.8842460, 0.1306200, 0.3485000, 0.3110900, 0.8564650, 0.7154170, 0.3940250, 0.7276840, 0.7968730, 0.7591330, 0.0364611, 0.3133540, 0.6116540, 0.1252610, 0.4822220, 0.1197930, 0.4094650, 0.4694960, 0.4545230, 0.2205010, 0.0755253, 0.9767120, 0.9914310, 0.0459867, 0.5205610, 0.0153277, 0.7233090, 0.7525990, 0.8137740, 0.8881650, 0.2331970, 0.3007880, 0.4838210, 0.6410550, 0.9055880, 0.2437180, 0.2624710, 0.2655750, 0.4483450, 0.7951410, 0.2621020, 0.8165700, 0.6718280, 0.6483310, 0.3906660, 0.4837060, 0.3457100, 0.9913590, 0.1446340, 0.6451250, 0.9062120, 0.9530850, 0.8012900, 0.8618790, 0.0488761, 0.9793320, 0.4424000, 0.5272520, 0.3068100, 0.4899010, 0.4657010, 0.4957290, 0.6549910, 0.6757360, 0.9947430, 0.6027150, 0.3960950, 0.9782550, 0.6975410, 0.9763810, 0.0434605, 0.4454890, 0.1019620, 0.6754800, 0.3445950, 0.7300180, 0.5931300, 0.2883430, 0.6517590, 0.1371680, 0.6399940, 0.4545100, 0.2650550, 0.9733320, 0.2690060, 0.4927860, 0.1526150, 0.3531390, 0.5717430, 0.2415940, 0.5051480, 0.5557870, 0.2619850, 0.3017210, 0.9336360, 0.0963557, 0.4634380, 0.8862740, 0.7134650, 0.9216480, 0.3522220, 0.2244210, 0.5971100, 0.7110200, 0.1104760, 0.0934760, 0.5407450, 0.8947490, 0.8209010, 0.9519340, 0.4973500, 0.1299500, 0.0944263, 0.1009230, 0.0599226, 0.8893270, 0.9442270, 0.1185050, 0.9643430, 0.5264980, 0.6445720, 0.9897940, 0.9976700, 0.8576110, 0.0836504, 0.6970720, 0.4859920, 0.0062545, 0.7394890, 0.2811470, 0.9250900, 0.8698560, 0.9329960, 0.9495160, 0.9229440, 0.8961780, 0.7744740, 0.7186700, 0.9109290, 0.8391840, 0.1881800, 0.2419840, 0.9675970, 0.1173670, 0.1492710, 0.0245217, 0.5216850, 0.0929769, 0.4828830, 0.0893908, 0.4824910, 0.3810410, 0.0940524, 0.9688800, 0.1303880, 0.9845220, 0.4427940, 0.3019080, 0.5652950, 0.9761590, 0.2622250, 0.8814410, 0.3949000, 0.6632340, 0.2840690, 0.4970430, 0.6699180, 0.2947030, 0.6886090, 0.0442514, 0.7109510, 0.6419550, 0.0406738, 0.0736680, 0.9311580, 0.7707480, 0.2244920, 0.3180100, 0.3275550, 0.9777840, 0.6036990, 0.1281990, 0.4515270, 0.9489680, 0.6739450, 0.7214510, 0.6005040, 0.8441940, 0.5858170, 0.7471430, 0.2760020, 0.7298190, 0.1907070, 0.4593850, 0.8045970, 0.6798990, 0.2601070, 0.0126904, 0.6731910, 0.9815910, 0.1180470, 0.4193760, 0.1576620, 0.7753870, 0.9497600, 0.8256110, 0.6033770, 0.1515860, 0.8153380, 0.9371540, 0.1850520, 0.3232410, 0.3853880, 0.4231760, 0.3597800, 0.0678210, 0.6735670, 0.4970500, 0.5768620, 0.2070500, 0.3426430, 0.0390466, 0.4897910, 0.5991540, 0.7133170, 0.1677030, 0.4193450, 0.1026510, 0.2999570, 0.9712850, 0.8907510, 0.9462940, 0.7714920, 0.8167580, 0.6441910, 0.0385524, 0.3140910, 0.5201140, 0.0462578, 0.7092260, 0.5536750, 0.9299590, 0.5944450, 0.7175690, 0.8534450, 0.2899460, 0.1684510, 0.3417640, 0.4746770, 0.0636942, 0.7177840, 0.4831020, 0.7369160, 0.8461440, 0.1957450, 0.1571110, 0.3830620, 0.4376010, 0.2187870, 0.8459670, 0.3968370, 0.7579590, 0.8326590, 0.1012120, 0.7063700, 0.3311260, 0.9431650, 0.9272640, 0.6544380, 0.1066640, 0.9044260, 0.6200150, 0.6324330, 0.8397850, 0.3245450, 0.0027007, 0.1561200, 0.5856590, 0.9769720, 0.1723810, 0.5450610, 0.1360080, 0.8935640, 0.4150230, 0.0607805, 0.3270310, 0.5735750, 0.8203480, 0.9603120, 0.3533360, 0.4234270, 0.0569615, 0.4651450, 0.0682401, 0.8263880, 0.8378220, 0.8807010, 0.5063950, 0.7247010, 0.7291140, 0.1829210, 0.1113620, 0.0584858, 0.5787680, 0.9755870, 0.1071750, 0.2147040, 0.0296183, 0.8319660, 0.7459730, 0.0535969, 0.3538030, 0.5367530, 0.7282110, 0.3712670, 0.7196420, 0.5555670, 0.4314280, 0.5301640, 0.8442260, 0.3965770, 0.8530560, 0.8749430, 0.1909930, 0.6940000, 0.0499580, 0.1260890, 0.3292400, 0.9339280, 0.3118520, 0.6462800, 0.5837600, 0.2932200, 0.1238640, 0.4793820, 0.1496250, 0.6781960, 0.1697440, 0.5858120, 0.4710320, 0.3128360, 0.1110760, 0.7676590, 0.9387090, 0.5023260, 0.3343780, 0.7775020, 0.5773320, 0.3871660, 0.3286580, 0.5691640, 0.3563510, 0.8356560, 0.4801370, 0.3884310, 0.9267070, 0.8451780, 0.4828190, 0.5323520, 0.1775700, 0.0376971, 0.6012840, 0.2827140, 0.9352990, 0.3844350, 0.9696150, 0.1483230, 0.1471850, 0.0426928, 0.4959290, 0.2372570, 0.8537700, 0.9776960, 0.3920940, 0.0847186, 0.7211570, 0.1864130, 0.0847904, 0.7422170, 0.6757520, 0.5756260, 0.9864830, 0.9754010, 0.4916960, 0.6151670, 0.3665300, 0.4714510, 0.0921263, 0.9858840, 0.6046540, 0.9839510, 0.4631040, 0.9522510, 0.2708670, 0.5404710, 0.5254930, 0.3305600, 0.5315350, 0.0556472, 0.5603850, 0.3159520, 0.7565710, 0.9188300, 0.0616884, 0.4410410, 0.4749030, 0.3459300, 0.7259080, 0.0544611, 0.1691150, 0.6489750, 0.0556556, 0.5492900, 0.0397673, 0.5257110, 0.7119000, 0.2527000, 0.7944310, 0.2391860, 0.6852790, 0.1850620, 0.5000260, 0.5416650, 0.7699000, 0.4680520, 0.1766200, 0.7330770, 0.1988380, 0.7726020, 0.7660260, 0.4651440, 0.6907970, 0.9061660, 0.1118100, 0.3690240, 0.6993030, 0.0576149, 0.9888900, 0.3043090, 0.2190210, 0.3429300, 0.0317769, 0.2039150, 0.6251810, 0.8538720, 0.7781390, 0.6497900, 0.1885250, 0.8870240, 0.8622050, 0.2672620, 0.3828960, 0.1036760, 0.1635530, 0.4936040, 0.2143460, 0.3461540, 0.1849680, 0.3839620, 0.6951800, 0.5665830, 0.9365000, 0.2242830, 0.7629470, 0.4568770, 0.0122766, 0.3188430, 0.7591250, 0.2944680, 0.0876849, 0.6158760, 0.4554200, 0.4708670, 0.7193540, 0.9626220, 0.1904770, 0.8165150, 0.6737510, 0.6988590, 0.5339760, 0.1992670, 0.6678050, 0.5093100, 0.2713240, 0.7776910, 0.9325290, 0.4492160, 0.8249680, 0.2549080, 0.2137210, 0.8881960, 0.5380550, 0.1116390, 0.2900170, 0.5964870, 0.1792680, 0.9172370, 0.6976610, 0.1722550, 0.8023020, 0.3920280, 0.0037012, 0.6575040, 0.8113920, 0.2654090, 0.2658660, 0.0761886, 0.4009630, 0.4584270, 0.8309220, 0.5977560, 0.1259870, 0.3978380, 0.9242490, 0.4869080, 0.7878220, 0.6490020, 0.0430807, 0.9086940, 0.1274720, 0.7205040, 0.4321060, 0.6872350, 0.9664940, 0.3949960, 0.8137770, 0.2891850, 0.5481450, 0.5621100, 0.9946710, 0.6886480, 0.3095230, 0.1298340, 0.8664830, 0.1004500, 0.8008420, 0.7034650, 0.3675800, 0.5135790, 0.2484130, 0.6620580, 0.9167580, 0.6445920, 0.8450620, 0.0411495, 0.6298600, 0.8996970, 0.1865210, 0.3324090, 0.0680878, 0.2073380, 0.6473490, 0.2095920, 0.5538880, 0.5878080, 0.0431148, 0.3812860, 0.5894030, 0.8448290, 0.1247340, 0.4192710, 0.8650400, 0.6984610, 0.9479950, 0.7586420, 0.5371630, 0.9723540, 0.3877120, 0.1904790, 0.2067200, 0.9438570, 0.1407760, 0.7576830, 0.3938260, 0.4222260, 0.4909350, 0.8787110, 0.8183690, 0.4058540, 0.1446670, 0.9513870, 0.9264710, 0.8668980, 0.9034370, 0.0897642, 0.0628556, 0.9153340, 0.9349180, 0.3514390, 0.8356020, 0.4851460, 0.1450950, 0.0976653, 0.5688510, 0.7470980, 0.1940000, 0.6207130, 0.1379970, 0.8006970, 0.9084410, 0.3323550, 0.1707720, 0.3303540, 0.8547460, 0.8688980, 0.7403530, 0.7378440, 0.7695770, 0.2780480, 0.9511920, 0.6427110, 0.5845110, 0.0466777, 0.1314160, 0.7127980, 0.4517230, 0.9600710, 0.3188980, 0.3135070, 0.3362330, 0.5349130, 0.1361860, 0.3682540, 0.5065310, 0.2837180, 0.4125180, 0.9058580, 0.3295960, 0.2127400, 0.5759330, 0.0461932, 0.0835102, 0.3423990, 0.7684190, 0.2205630, 0.1451710, 0.8833790, 0.1923550, 0.8287690, 0.8158520, 0.1347670, 0.0625876, 0.6750830, 0.5353660, 0.4465640, 0.0810434, 0.9996070, 0.1006660, 0.0384967, 0.3188980, 0.0775650, 0.3846520, 0.1118410, 0.9324660, 0.3335360, 0.9986240, 0.3490520, 0.6644580, 0.1979980, 0.5048130, 0.3395830, 0.7581720, 0.5890200, 0.2090200, 0.1582680, 0.9179290, 0.3220950, 0.3910110, 0.5860440, 0.4732530, 0.4485400, 0.5071690, 0.7583270, 0.9665040, 0.6990900, 0.6361660, 0.7629190, 0.0959780, 0.9250400, 0.3141480, 0.0427695, 0.1054420, 0.4182410, 0.4820330, 0.4107140, 0.3398060, 0.3113430, 0.5966920, 0.1184920, 0.7111080, 0.5555070, 0.3374270, 0.6907840, 0.9805960, 0.9794310, 0.5998390, 0.7405270, 0.4858850, 0.2624090, 0.5592240, 0.8890640, 0.1893230, 0.2810180, 0.8053880, 0.3876100, 0.3748390, 0.5092730, 0.4320050, 0.2467080, 0.0652057, 0.1061540, 0.3227290, 0.8348730, 0.3703290, 0.9074230, 0.2190920, 0.6273990, 0.4448100, 0.8098460, 0.5917280, 0.9617850, 0.9641880, 0.6727580, 0.1290390, 0.3751820, 0.2331720, 0.4963960, 0.9937830, 0.7772210, 0.1998260, 0.8513000, 0.8086100, 0.9539270, 0.3052140, 0.4079300, 0.6733840, 0.5672080, 0.7222220, 0.7309600, 0.1581200, 0.0427850, 0.7623220, 0.5271890, 0.8421310, 0.7210180, 0.2663280, 0.7928500, 0.3413980, 0.6704540, 0.3514690, 0.8795780, 0.0192828, 0.3092920, 0.0492666, 0.2022930, 0.8626340, 0.7779490, 0.0455279, 0.4162000, 0.7271130, 0.9194360, 0.4204900, 0.1582370, 0.7575210, 0.4919290, 0.1381920, 0.1978130, 0.9298010, 0.8847910, 0.7100220, 0.6682310, 0.4189010, 0.2674120, 0.3869220, 0.7132320, 0.7152710, 0.5478640, 0.5945730, 0.7431310, 0.6076240, 0.2263120, 0.0328178, 0.6179280, 0.6385360, 0.1552320, 0.2825290, 0.1260240, 0.3504870, 0.5214060, 0.0342883, 0.2939340, 0.8253880, 0.5987110, 0.8607230, 0.7495990, 0.1889770, 0.0965978, 0.6221940, 0.0458032, 0.1132730, 0.0803912, 0.9328780, 0.5058820, 0.3652970, 0.2537630, 0.9811690, 0.0077981, 0.9543570, 0.7995680, 0.1937610, 0.9169540, 0.3357710, 0.1358260, 0.7967540, 0.3826940, 0.9219750, 0.6423780, 0.6972770, 0.0120370, 0.2385000, 0.9468390, 0.0894302, 0.7006670, 0.5991610, 0.2755720, 0.1262300, 0.4116590, 0.1344580, 0.1348520, 0.3998330, 0.3653540, 0.8621060, 0.6029790, 0.1525210, 0.0205639, 0.8161680, 0.5281990, 0.9571170, 0.8234250, 0.4418740, 0.5425150, 0.5958320, 0.4175780, 0.3495680, 0.1490360, 0.0881526, 0.4283380, 0.0417103, 0.6528980, 0.2622980, 0.0899725, 0.7679490, 0.1883430, 0.4577670, 0.7424010, 0.1813170, 0.3716260, 0.7116830, 0.5133040, 0.9817440, 0.6987230, 0.1189870, 0.5337560, 0.6096360, 0.9973210, 0.8364430, 0.7751330, 0.8867220, 0.9109290, 0.0587728, 0.0997106, 0.1504600, 0.5932370, 0.2602540, 0.6445910, 0.6970780, 0.5322130, 0.5650010, 0.7879130, 0.9620280, 0.8604190, 0.4501660, 0.1940940, 0.9274310, 0.5491040, 0.4048070, 0.4249270, 0.5648730, 0.7935010, 0.6842290, 0.0208552, 0.0478051, 0.8074330, 0.3847780, 0.4618040, 0.1783560, 0.2782910, 0.0668262, 0.5873710, 0.2508250, 0.3204120, 0.8486270, 0.3218400, 0.8489410, 0.5656770, 0.9310230, 0.3683670, 0.0211677, 0.7583570, 0.8813600, 0.6318190, 0.9833680, 0.3720780, 0.8962820, 0.7752270, 0.1818790, 0.2160160, 0.1805770, 0.3651250, 0.4110410, 0.4461780, 0.1140010, 0.7712140, 0.7684640, 0.7503030, 0.7529630, 0.7266540, 0.5393480, 0.3722660, 0.9905100, 0.7620950, 0.0047922, 0.6933260, 0.4743310, 0.1678070, 0.0483881, 0.2253510, 0.7655190, 0.0889216, 0.2519360, 0.9013820, 0.3881090, 0.0925243, 0.7070760, 0.1298250, 0.2749590, 0.1998890, 0.2759100, 0.8759690, 0.5586280, 0.8893790, 0.3012710, 0.8941490, 0.6976130, 0.7043470, 0.1088890, 0.4157830, 0.6891730, 0.4763700, 0.3878210, 0.4071130, 0.4897500, 0.1858650, 0.1040310, 0.5760770, 0.8851690, 0.2044910, 0.5349960, 0.5476150, 0.3633290, 0.6405170, 0.3211070, 0.0335866, 0.3257970, 0.8356450, 0.1927340, 0.6442890, 0.9685100, 0.6952700, 0.5725180, 0.5908020, 0.2685890, 0.0474654, 0.8558730, 0.5692040, 0.6883660, 0.9572140, 0.6867850, 0.0007137, 0.9096650, 0.8973330, 0.8240700, 0.4056330, 0.5911020, 0.2984200, 0.7811230, 0.6897000, 0.9358740, 0.2358730, 0.9838590, 0.4143400, 0.9799110, 0.0791655, 0.0578072, 0.5441010, 0.3987900, 0.6455640, 0.6870700, 0.0891235, 0.4661920, 0.4199950, 0.0649898, 0.3680590, 0.3003300, 0.7674390, 0.1057500, 0.6375020, 0.8548240, 0.2401890, 0.6560260, 0.5609040, 0.9331600, 0.1392720, 0.8765580, 0.3811730, 0.3831030, 0.3185560, 0.2535560, 0.2152630, 0.9547860, 0.1600510, 0.4579860, 0.1284310, 0.2057920, 0.3988790, 0.3083800, 0.7911710, 0.9600650, 0.5256000, 0.5303940, 0.8615830, 0.0521196, 0.1239040, 0.9099380, 0.9464000, 0.9681020, 0.4968190, 0.3449360, 0.3506400, 0.0215136, 0.5080490, 0.5428000, 0.7306120, 0.9130610, 0.6400020, 0.8206450, 0.5436700, 0.5755450, 0.7334500, 0.0975657, 0.4442050, 0.9409920, 0.0215130, 0.5939040, 0.2779970, 0.8464100, 0.4704590, 0.1666410, 0.5087130, 0.7932800, 0.4814850, 0.8871470, 0.4007150, 0.3590220, 0.5036150, 0.9512880, 0.0794576, 0.5106700, 0.0134271, 0.7935780, 0.3610910, 0.9936140, 0.0200632, 0.5677210, 0.1610550, 0.7897830, 0.9610630, 0.4104350, 0.1711600, 0.2620340, 0.4945230, 0.1600580, 0.5075630, 0.1539520, 0.1696490, 0.2949830, 0.9381970, 0.2816110, 0.1183780, 0.7098190, 0.0421854, 0.5818710, 0.5296480, 0.5842370, 0.6827700, 0.8951670, 0.7856330, 0.4372500, 0.7265340, 0.5093950, 0.8381860, 0.3829550, 0.4801060, 0.8690590, 0.4956310, 0.6089820, 0.6492110, 0.0202991, 0.7592260, 0.9056730, 0.1569470, 0.5128230, 0.7616660, 0.0152500, 0.2900460, 0.9193100, 0.5130870, 0.0284486, 0.0404045, 0.2253670, 0.2518490, 0.1315280, 0.7525490, 0.3201860, 0.4180300, 0.8192460, 0.1187990, 0.1663470, 0.8239390, 0.1900420, 0.1936840, 0.6432920, 0.6008590, 0.5922400, 0.5896560, 0.3930390, 0.3798280, 0.9110000, 0.4736370, 0.3921500, 0.3467060, 0.9077310, 0.3129040, 0.5191380, 0.9740950, 0.4740320, 0.6175610, 0.1710750, 0.9289060, 0.4065080, 0.1148660, 0.8056320, 0.0207510, 0.1296420, 0.2165430, 0.6926650, 0.8081420, 0.2938060, 0.4740710, 0.5798710, 0.6105430, 0.0912483, 0.2681460, 0.8492210, 0.4707640, 0.2898650, 0.3023900, 0.8703670, 0.4807090, 0.6843190, 0.9582900, 0.8122280, 0.3300320, 0.3894800, 0.1765880, 0.3324710, 0.7354120, 0.0157217, 0.0853309, 0.1976220, 0.8409720, 0.3209250, 0.3598290, 0.2201710, 0.7433090, 0.1543230, 0.1289140, 0.3204500, 0.2865820, 0.0483622, 0.3391080, 0.4742460, 0.1784690, 0.9963780, 0.2362170, 0.5617660, 0.8430010, 0.3472150, 0.3055980, 0.9848000, 0.1198130, 0.2567540, 0.0498737, 0.2277520, 0.2796250, 0.3155990, 0.9783760, 0.0859696, 0.6490060, 0.1672100, 0.6761070, 0.7847970, 0.2997610, 0.6447930, 0.0538474, 0.4515170, 0.2386240, 0.6432930, 0.6719670, 0.7413000, 0.3483260, 0.0741213, 0.9939900, 0.9189460, 0.2204410, 0.1428380, 0.5584380, 0.7249420, 0.1217220, 0.5194780, 0.0869088, 0.6376140, 0.4395930, 0.9682090, 0.7552030, 0.6295950, 0.1851770, 0.1378810, 0.6657740, 0.4027190, 0.5136770, 0.8671570, 0.4573140, 0.0438009, 0.0773345, 0.8289830, 0.0375343, 0.4013120, 0.1533890, 0.7631410, 0.6667250, 0.0682487, 0.3160270, 0.4774800, 0.8916880, 0.7343780, 0.4473140, 0.7625530, 0.7391490, 0.1222640, 0.4055080, 0.5245200, 0.5534560, 0.4982430, 0.1372870, 0.1152460, 0.8657620, 0.4113820, 0.3972270, 0.5696680, 0.0987829, 0.5738690, 0.6878870, 0.5725980, 0.3953270, 0.4643000, 0.8629910, 0.6683550, 0.4113600, 0.7454440, 0.7554060, 0.4809370, 0.1344670, 0.2897940, 0.8551540, 0.7452700, 0.0352387, 0.1643480, 0.2754490, 0.2321170, 0.1578880, 0.6739800, 0.9084800, 0.7708190, 0.8004940, 0.9927480, 0.9105130, 0.9485460, 0.5104630, 0.8025170, 0.5735220, 0.8660810, 0.8365520, 0.6954390, 0.8434810, 0.3673860, 0.5211880, 0.3943550, 0.4409410, 0.7810350, 0.0498857, 0.0489585, 0.5611210, 0.2050500, 0.8438120, 0.1842800, 0.5760050, 0.2410530, 0.3115750, 0.9293160, 0.1692480, 0.7138940, 0.5771830, 0.6126190, 0.9677710, 0.3164160, 0.1644120, 0.4057920, 0.5441850, 0.4005760, 0.3604600, 0.9549040, 0.2503560, 0.8046010, 0.7367510, 0.7179690, 0.0635708, 0.0073857, 0.1562500, 0.9590330, 0.9141260, 0.3073320, 0.1961500, 0.1812420, 0.5290270, 0.5735840, 0.7944250, 0.9306260, 0.9060210, 0.7888330, 0.1294380, 0.2096640, 0.8957200, 0.6675360, 0.6372570, 0.6028650, 0.1539260, 0.8744400, 0.5718500, 0.7933160, 0.4249050, 0.3951370, 0.4103930, 0.6596270, 0.0630654, 0.0591461, 0.6004390, 0.0954817, 0.3600590, 0.8696470, 0.8302870, 0.3591180, 0.9298490, 0.7068090, 0.7322070, 0.5249100, 0.9411580, 0.4818930, 0.5092560, 0.5897240, 0.3825150, 0.6522690, 0.9106290, 0.0522056, 0.7902810, 0.8888290, 0.0152475, 0.0457682, 0.4479800, 0.8330720, 0.2916950, 0.8757160, 0.3113340, 0.4381680, 0.5526010, 0.7402680, 0.8118750, 0.1869420, 0.7508740, 0.2312270, 0.0601643, 0.3306880, 0.3933270, 0.6657360, 0.2646580, 0.0707114, 0.9244370, 0.3816660, 0.3954710, 0.2646880, 0.7309430, 0.1047340, 0.0636853, 0.2205760, 0.4632770, 0.4969420, 0.5268380, 0.1033350, 0.8818730, 0.1973420, 0.2305160, 0.4871090, 0.0230257, 0.9665780, 0.1956070, 0.9626670, 0.8859460, 0.6910160, 0.5265680, 0.4115980, 0.0265164, 0.6777750, 0.5798690, 0.4908850, 0.9876300, 0.3101600, 0.9986050, 0.8796260, 0.3617620, 0.2277120, 0.6984450, 0.1825180, 0.7145320, 0.1066950, 0.5645090, 0.7054060, 0.4936350, 0.2714030, 0.9613490, 0.9861090, 0.2584090, 0.2272750, 0.1848470, 0.2578840, 0.9813780, 0.4949740, 0.5169680, 0.2947580, 0.1787300, 0.7964360, 0.9938890, 0.0187124, 0.8785430, 0.4570140, 0.5211500, 0.6593040, 0.9316170, 0.8802270, 0.2321610, 0.7644710, 0.6603980, 0.4871340, 0.4038320, 0.3157910, 0.0616432, 0.1669490, 0.9146720, 0.2288610, 0.6677100, 0.3045690, 0.0214811, 0.6680960, 0.2113140, 0.9572140, 0.5641310, 0.1141500, 0.5435800, 0.1258800, 0.3502730, 0.1922060, 0.4623020, 0.5409440, 0.0039512, 0.9647720, 0.5028330, 0.5861110, 0.9696830, 0.8362980, 0.5920570, 0.5786880, 0.0494181, 0.6472230, 0.6319530, 0.0654165, 0.7789150, 0.0228701, 0.6582190, 0.2747820, 0.3901070, 0.6809710, 0.0018287, 0.2713840, 0.2019520, 0.1026160, 0.4410410, 0.8781110, 0.2242450, 0.6498480, 0.3456640, 0.9533640, 0.7428260, 0.5607760, 0.1848250, 0.8472850, 0.1088760, 0.3714590, 0.4113260, 0.7902000, 0.4594590, 0.1332830, 0.4864180, 0.3132250, 0.7779660, 0.1735420, 0.8633820, 0.7702140, 0.3111700, 0.4771720, 0.9686220, 0.6377230, 0.8349560, 0.3501600, 0.3141500, 0.9782010, 0.3095570, 0.9763570, 0.5690060, 0.4887810, 0.5299210, 0.7934740, 0.4596750, 0.1347550, 0.9463390, 0.1292780, 0.6355550, 0.0648678, 0.8677510, 0.3976790, 0.6961170, 0.0849685, 0.8039750, 0.1123760, 0.9734020, 0.9975780, 0.0399340, 0.5379130, 0.0252336, 0.1742110, 0.9302400, 0.0280736, 0.5404350, 0.3107210, 0.7488160, 0.1498740, 0.1908100, 0.4484370, 0.1673570, 0.3125870, 0.9327720, 0.4656890, 0.4485860, 0.4008810, 0.5763940, 0.0790341, 0.5559170, 0.7884370, 0.3824060, 0.0228641, 0.5978680, 0.0354778, 0.8841210, 0.0391017, 0.7833920, 0.4624710, 0.3475840, 0.9438230, 0.9516110, 0.7140940, 0.5964810, 0.7697140, 0.9773360, 0.2687300, 0.4057280, 0.8289990, 0.2697410, 0.0026182, 0.4357570, 0.4257050, 0.2133140, 0.2472700, 0.5136300, 0.9508410, 0.5779730, 0.5746150, 0.4167400, 0.2154170, 0.7012890, 0.5813750, 0.0785233, 0.0986814, 0.7729080, 0.1402020, 0.4679310, 0.4815270, 0.1645460, 0.5701830, 0.1762380, 0.0930225, 0.8040390, 0.2992150, 0.2920220, 0.1753530, 0.0412818, 0.7877870, 0.5670960, 0.2933310, 0.0474824, 0.3225760, 0.0661163, 0.6674330, 0.4625880, 0.2505000, 0.9230920, 0.3384590, 0.9976380, 0.4868600, 0.6237620, 0.9110770, 0.1275090, 0.2864320, 0.9004950, 0.8545920, 0.7326070, 0.1397100, 0.1635420, 0.4828840, 0.2166380, 0.2492610, 0.3234250, 0.3554520, 0.6054990, 0.8185720, 0.5869140, 0.1908380, 0.3465030, 0.7880990, 0.2239430, 0.9013490, 0.0349908, 0.1864680, 0.7956930, 0.4663070, 0.2000200, 0.5692550, 0.0088515, 0.2355070, 0.3244070, 0.4118940, 0.2684730, 0.3496470, 0.9636450, 0.3941960, 0.4085180, 0.5599010, 0.5668200, 0.4696400, 0.3506420, 0.5322650, 0.7877090, 0.4812750, 0.7036110, 0.7554780, 0.0857419, 0.8703800, 0.6209170, 0.8732090, 0.2157820, 0.5412900, 0.6161220, 0.2945380, 0.7707060, 0.9547420, 0.9385410, 0.3016670, 0.4264550, 0.5749580, 0.1617080, 0.9128490, 0.2069260, 0.5914830, 0.1601480, 0.2865050, 0.4748470, 0.4350780, 0.7999390, 0.7580650, 0.4022880, 0.4543210, 0.4762280, 0.9014440, 0.9695660, 0.5229590, 0.0699167, 0.3750540, 0.3588610, 0.2023680, 0.0097718, 0.8815680, 0.6100340, 0.2485730, 0.7218600, 0.8606660, 0.2501730, 0.9295410, 0.6191930, 0.0263395, 0.4358280, 0.2556770, 0.0749437, 0.4805910, 0.7404580, 0.9144790, 0.4751540, 0.7926550, 0.7687380, 0.7956860, 0.3118730, 0.0768719, 0.5503540, 0.2278290, 0.5461730, 0.2357480, 0.4894830, 0.1480700, 0.2258930, 0.8531280, 0.2349700, 0.5281060, 0.7848460, 0.5815220, 0.9160060, 0.8863310, 0.1931680, 0.9466820, 0.1461860, 0.9037350, 0.1643400, 0.4368330, 0.2253510, 0.6594740, 0.6524750, 0.3240900, 0.7872660, 0.1683430, 0.0174890, 0.6904800, 0.8440340, 0.3162610, 0.9261170, 0.6421520, 0.3928480, 0.6696870, 0.9254620, 0.9757540, 0.1013350, 0.4108300, 0.5675280, 0.0986873, 0.4525960, 0.6343200, 0.3840660, 0.2024330, 0.7083290, 0.1469970, 0.2493150, 0.9904530, 0.4894370, 0.8183370, 0.3304220, 0.3196100, 0.2491510, 0.3216930, 0.3872010, 0.5074420, 0.0180923, 0.0548384, 0.8912890, 0.7260440, 0.2437930, 0.1236130, 0.1246770, 0.9365050, 0.3562450, 0.5088020, 0.4348430, 0.1256750, 0.5242360, 0.3364770, 0.9990540, 0.0385927, 0.9139900, 0.0712975, 0.2666140, 0.9529210, 0.0559188, 0.6475460, 0.2824350, 0.5695030, 0.9271900, 0.4877500, 0.8793530, 0.0338833, 0.7651090, 0.5394930, 0.5158330, 0.7458220, 0.3923320, 0.9520390, 0.8608700, 0.9010980, 0.7168860, 0.3839740, 0.2739100, 0.6369560, 0.2714710, 0.4464280, 0.4828250, 0.5722800, 0.5281300, 0.8301440, 0.2282820, 0.4237770, 0.6163050, 0.4296360, 0.2711910, 0.1428290, 0.9727820, 0.0775685, 0.1501110, 0.3506980, 0.3440330, 0.5371930, 0.1661830, 0.3758090, 0.4519180, 0.7639880, 0.7779670, 0.2831150, 0.9379920, 0.7471120, 0.2203920, 0.8020510, 0.7404450, 0.3980270, 0.1811070, 0.1500620, 0.9167290, 0.7592640, 0.9035240, 0.7269620, 0.6953360, 0.4612770, 0.8034800, 0.4315070, 0.0450203, 0.6367390, 0.5141000, 0.7934030, 0.2357400, 0.2354230, 0.7235250, 0.0721295, 0.7781050, 0.6141490, 0.5712070, 0.6670250, 0.8316730, 0.2522610, 0.7022880, 0.8334520, 0.6777340, 0.6709490, 0.6717350, 0.1398780, 0.2035500, 0.9644750, 0.1733440, 0.4480410, 0.5988310, 0.5865230, 0.0183551, 0.2049030, 0.2155880, 0.1960360, 0.2154900, 0.5114450, 0.4621280, 0.0446196, 0.5387420, 0.9705780, 0.2207940, 0.5708400, 0.9403000, 0.3792040, 0.7524500, 0.4998940, 0.7735780, 0.3515110, 0.7164100, 0.1649580, 0.5968650, 0.7430420, 0.8337710, 0.9958010, 0.9940930, 0.0813356, 0.1728560, 0.6698460, 0.2517870, 0.5963380, 0.5456860, 0.9013490, 0.9945630, 0.9783110, 0.4505300, 0.5412400, 0.8729020, 0.9821070, 0.6223230, 0.6355190, 0.6772710, 0.4105440, 0.7683760, 0.5030640, 0.2033800, 0.7423890, 0.8270990, 0.4048740, 0.8993450, 0.8775700, 0.9074810, 0.1741580, 0.1984590, 0.5028400, 0.0332960, 0.8782370, 0.3090650, 0.7242080, 0.2067850, 0.2842100, 0.3125180, 0.9770670, 0.4823500, 0.6273230, 0.3711560, 0.6911010, 0.0376874, 0.1916940, 0.0913877, 0.6654130, 0.6052830, 0.8853000, 0.0420876, 0.6528380, 0.3248510, 0.2463940, 0.4497330, 0.7859690, 0.8617340, 0.5155540, 0.8182430, 0.7026710, 0.9816740, 0.6805340, 0.6494370, 0.3556010, 0.5139850, 0.0740471, 0.7423260, 0.8596820, 0.6748730, 0.2674680, 0.1648820, 0.4126960, 0.2386380, 0.3982580, 0.3039860, 0.1777350, 0.9481750, 0.8164000, 0.5523160, 0.9240390, 0.3959830, 0.2051620, 0.2131290, 0.5159880, 0.7595630, 0.6562310, 0.1721640, 0.6144030, 0.4752100, 0.1741610, 0.4415530, 0.3535710, 0.3825970, 0.5137770, 0.9700350, 0.3586400, 0.5629240, 0.8079360, 0.6236850, 0.1995550, 0.4538810, 0.9181450, 0.7687580, 0.9224160, 0.3916040, 0.9788760, 0.9869220, 0.4430250, 0.1339530, 0.5121400, 0.3028120, 0.5292970, 0.4883240, 0.6903930, 0.5733440, 0.0779331, 0.7132670, 0.0839810, 0.1121820, 0.3494450, 0.2512430, 0.5048560, 0.2001900, 0.5734450, 0.4927270, 0.2240100, 0.3595830, 0.2520470, 0.4084060, 0.2639070, 0.9994810, 0.1740130, 0.9374150, 0.0109464, 0.2124690, 0.3055840, 0.8997730, 0.9309900, 0.4507770, 0.0998693, 0.9249710, 0.2874870, 0.1079480, 0.6446440, 0.8813970, 0.1502380, 0.7078460, 0.6468080, 0.0009778, 0.2417720, 0.2044470, 0.0836219, 0.2035000, 0.7251050, 0.3489480, 0.0049560, 0.6328920, 0.2966500, 0.6619390, 0.1043180, 0.0657007, 0.2758610, 0.3483250, 0.1002960, 0.7433060, 0.8900320, 0.0857892, 0.5659320, 0.0963086, 0.8757930, 0.4595020, 0.4540590, 0.1083600, 0.0296070, 0.2189090, 0.5415020, 0.9456410, 0.5836690, 0.1960630, 0.3432300, 0.8187340, 0.3786610, 0.4968890, 0.7656780, 0.5304030, 0.2440220, 0.4287530, 0.1485560, 0.4533430, 0.0612332, 0.1055260, 0.1775990, 0.7454550, 0.4656130, 0.0901638, 0.7880370, 0.8157640, 0.6872140, 0.7264890, 0.3141530, 0.6293430, 0.3929360, 0.7297240, 0.7273670, 0.1039120, 0.5685400, 0.0626407, 0.4473230, 0.5706750, 0.5734700, 0.7802560, 0.2619850, 0.2810130, 0.0035031, 0.4334950, 0.8712440, 0.7617870, 0.7023300, 0.1037150, 0.8462200, 0.2527910, 0.1375990, 0.9066380, 0.8327340, 0.0820183, 0.2989910, 0.3761620, 0.0479592, 0.5408350, 0.1410500, 0.6955410, 0.0770796, 0.9458130, 0.1148230, 0.8229930, 0.5103240, 0.6427750, 0.3498660, 0.2965490, 0.3443490, 0.9093280, 0.2208950, 0.9095350, 0.4130930, 0.0428756, 0.2741470, 0.8103410, 0.7714570, 0.9318410, 0.3384820, 0.8422500, 0.3875300, 0.5206030, 0.3646500, 0.5597450, 0.2941940, 0.2014130, 0.0211083, 0.9246680, 0.1082810, 0.0324374, 0.1771050, 0.8265530, 0.0765446, 0.1279820, 0.6574120, 0.4705400, 0.0202671, 0.5932480, 0.3405440, 0.2610030, 0.5975150, 0.0830871, 0.8331490, 0.5413460, 0.6248010, 0.8332490, 0.8089350, 0.2726500, 0.8199800, 0.3951860, 0.4209840, 0.3429550, 0.2460060, 0.7746330, 0.3505920, 0.8406480, 0.1358630, 0.4633700, 0.8559500, 0.4796990, 0.1239130, 0.7536690, 0.7293910, 0.8945600, 0.5218100, 0.7073380, 0.0262126, 0.3031970, 0.2417640, 0.8610900, 0.9260750, 0.2658060, 0.7359700, 0.1980990, 0.4493780, 0.3588000, 0.6465960, 0.7180170, 0.4222090, 0.8915490, 0.4007890, 0.7338120, 0.5199180, 0.5245250, 0.7235610, 0.8200120, 0.3664080, 0.3628630, 0.9471380, 0.8276740, 0.0344346, 0.9960380, 0.6236440, 0.1132420, 0.4953560, 0.3038310, 0.0814047, 0.4046200, 0.0680598, 0.9950490, 0.0586573, 0.1743080, 0.2027050, 0.5143460, 0.9404080, 0.1334240, 0.1376180, 0.5256430, 0.9620780, 0.8574920, 0.8600280, 0.7282700, 0.6988430, 0.9916900, 0.6051850, 0.5764750, 0.8114340, 0.8820780, 0.9850350, 0.5483080, 0.6478750, 0.2598890, 0.6069560, 0.6563260, 0.9397160, 0.1804400, 0.5682200, 0.7017260, 0.0914514, 0.6537880, 0.4503400, 0.5313760, 0.6825330, 0.7154620, 0.4006290, 0.1918410, 0.3759140, 0.9728460, 0.3411620, 0.2759520, 0.3112530, 0.0985604, 0.1369010, 0.3803280, 0.5321340, 0.2578570, 0.4746250, 0.9329140, 0.3463670, 0.3548910, 0.8197700, 0.1169620, 0.1465420, 0.8578730, 0.6147080, 0.2180050, 0.7977830, 0.3928550, 0.9972440, 0.7219110, 0.6957710, 0.1673620, 0.8337000, 0.5855470, 0.7608000, 0.3003280, 0.8639210, 0.6785100, 0.5382610, 0.5131760, 0.4541320, 0.8660280, 0.1983190, 0.6027010, 0.3963410, 0.6477340, 0.5641440, 0.8000310, 0.1812860, 0.6636350, 0.0493417, 0.0673879, 0.3250310, 0.5546960, 0.3548550, 0.6625650, 0.1449930, 0.5992220, 0.0241262, 0.8544320, 0.9512250, 0.1087570, 0.9451280, 0.8164610, 0.9521660, 0.3770330, 0.4668080, 0.9694670, 0.9707310, 0.2069050, 0.6878530, 0.1301310, 0.5678690, 0.1234740, 0.8561990, 0.0974818, 0.6246120, 0.7612030, 0.8717050, 0.3027540, 0.9954290, 0.4550940, 0.5382130, 0.9914360, 0.4818010, 0.2892550, 0.1151120, 0.8581040, 0.6431550, 0.7045920, 0.8515360, 0.3755740, 0.3851030, 0.1565460, 0.8939120, 0.1682440, 0.7423240, 0.5363900, 0.7524060, 0.2899830, 0.5257610, 0.8999180, 0.4222220, 0.9885140, 0.5243940, 0.2488650, 0.6079830, 0.0454191, 0.8303270, 0.1819830, 0.5667640, 0.9844430, 0.8909360, 0.8199980, 0.1938230, 0.4306660, 0.3510790, 0.8559790, 0.7433590, 0.8885870, 0.9016100, 0.2999680, 0.9083440, 0.4087430, 0.3586420, 0.2442980, 0.1314010, 0.1926080, 0.6754350, 0.7669390, 0.9637910, 0.5682360, 0.9515240, 0.6981530, 0.5053510, 0.5924850, 0.5781600, 0.6822980, 0.2758780, 0.5861730, 0.5359240, 0.0652490, 0.2885290, 0.1053420, 0.4398210, 0.3432240, 0.0384978, 0.2383810, 0.4821420, 0.6441740, 0.4858920, 0.5348260, 0.5352670, 0.0563633, 0.4060450, 0.2334830, 0.0402745, 0.2224910, 0.9536960, 0.9540970, 0.8468680, 0.3148920, 0.6940930, 0.6546160, 0.5035490, 0.4034170, 0.7708900, 0.0134790, 0.8833240, 0.3189010, 0.6576120, 0.5983860, 0.4057880, 0.4201530, 0.9725110, 0.4269590, 0.7726360, 0.8437930, 0.1171820, 0.8964660, 0.9868340, 0.0349061, 0.2331770, 0.2961670, 0.1714930, 0.0656071, 0.9102190, 0.6285390, 0.0892658, 0.8682830, 0.4691700, 0.0834424, 0.7165070, 0.0309399, 0.4709710, 0.7327930, 0.8592530, 0.5876750, 0.1125480, 0.7524180, 0.4801550, 0.5377360, 0.5809300, 0.7022340, 0.9290890, 0.3112650, 0.4015350, 0.6767960, 0.0275089, 0.9388070, 0.4501720, 0.8287960, 0.5765130, 0.8222490, 0.9760380, 0.0167127, 0.4758420, 0.2005640, 0.7094730, 0.1969750, 0.9557800, 0.3525470, 0.8419080, 0.9170050, 0.4430470, 0.5489190, 0.6424890, 0.9066030, 0.0940650, 0.9823600, 0.5524510, 0.5769490, 0.9468120, 0.9721010, 0.8800400, 0.0407743, 0.3969660, 0.8204580, 0.7042170, 0.9300920, 0.1473580, 0.6010870, 0.7345340, 0.1726090, 0.4306870, 0.9981720, 0.1323060, 0.5041810, 0.8469740, 0.8435190, 0.4733250, 0.8470860, 0.3067790, 0.3487180, 0.3753710, 0.5241010, 0.2349360, 0.8332820, 0.9685930, 0.6182680, 0.2297420, 0.9859390, 0.2848530, 0.0623202, 0.3152890, 0.7805510, 0.0408610, 0.5164310, 0.7061300, 0.2647960, 0.1597240, 0.7018330, 0.1117920, 0.9056130, 0.8015810, 0.2432780, 0.6196620, 0.0960803, 0.4424860, 0.0618646, 0.6223970, 0.2552120, 0.1781380, 0.7538720, 0.9335870, 0.9079360, 0.6436800, 0.6356280, 0.7674360, 0.6190830, 0.8978450, 0.1507520, 0.2404630, 0.8625540, 0.4378160, 0.4222640, 0.3886260, 0.7332400, 0.3409550, 0.8422290, 0.9110520, 0.5517100, 0.9327350, 0.2125730, 0.5671920, 0.1072810, 0.1568220, 0.1608610, 0.1659200, 0.7884290, 0.0808161, 0.5095400, 0.5639370, 0.2654060, 0.5917460, 0.5396710, 0.9402050, 0.4601890, 0.7243670, 0.1656780, 0.5029530, 0.3227630, 0.7595340, 0.6969790, 0.2404540, 0.9980480, 0.9084750, 0.3787620, 0.4423730, 0.0946736, 0.9216850, 0.0528245, 0.1042280, 0.1732470, 0.1181490, 0.0516227, 0.0535173, 0.4014940, 0.8136190, 0.8288870, 0.3327030, 0.0156800, 0.8533210, 0.5894470, 0.4920540, 0.1573600, 0.3531910, 0.9331170, 0.5418090, 0.7847220, 0.2405460, 0.4075620, 0.2544170, 0.2096490, 0.0085541, 0.1282170, 0.0683989, 0.2049270, 0.0678469, 0.4636590, 0.4746350, 0.4755270, 0.1806790, 0.3703050, 0.2597200, 0.1586740, 0.5121040, 0.5473850, 0.9875860, 0.3880020, 0.7556330, 0.4733300, 0.2679690, 0.9188590, 0.0279915, 0.5617710, 0.5865590, 0.2252610, 0.9081050, 0.6787980, 0.3566580, 0.5706620, 0.4263010, 0.6555830, 0.7592460, 0.5796620, 0.3940970, 0.1596040, 0.3477210, 0.5444660, 0.9773580, 0.4124280, 0.1823610, 0.0806040, 0.3641790, 0.8574120, 0.8683370, 0.3808830, 0.6678380, 0.4712060, 0.0148180, 0.8931800, 0.6960090, 0.5327030, 0.1902270, 0.0775560, 0.6480140, 0.9675050, 0.1838650, 0.6887260, 0.1249660, 0.1210610, 0.8984280, 0.6561990, 0.5042390, 0.1864610, 0.8091260, 0.5060780, 0.9872250, 0.3902490, 0.0745781, 0.4286450, 0.6432880, 0.7119790, 0.6438980, 0.3314740, 0.8041000, 0.2671320, 0.1110640, 0.9962840, 0.6407220, 0.5361970, 0.9683280, 0.3417850, 0.0558588, 0.2234850, 0.6605530, 0.8128160, 0.2901060, 0.8024860, 0.4449250, 0.1049200, 0.5298630, 0.4919430, 0.8144810, 0.7670050, 0.2056020, 0.2654750, 0.6786890, 0.3614590, 0.7052900, 0.2633440, 0.4461590, 0.2470630, 0.5606220, 0.2423010, 0.3848760, 0.9796950, 0.2911260, 0.8237020, 0.3158740, 0.2445890, 0.0198518, 0.6088170, 0.9820840, 0.1114240, 0.2235610, 0.6501550, 0.5242140, 0.7046600, 0.3709050, 0.7310390, 0.8502290, 0.0953953, 0.1517460, 0.9246320, 0.4000340, 0.4072300, 0.4105930, 0.2294270, 0.9370230, 0.1302670, 0.4552070, 0.7148800, 0.9915760, 0.1980560, 0.2757400, 0.6750800, 0.1873410, 0.0731626, 0.3862630, 0.2603130, 0.8070350, 0.5500810, 0.4474700, 0.3513260, 0.4581340, 0.4697390, 0.8566080, 0.1544500, 0.0451153, 0.7464510, 0.9527390, 0.7381840, 0.3096000, 0.7665420, 0.8041050, 0.9085610, 0.0691179, 0.9029200, 0.6281020, 0.5191220, 0.4902810, 0.3909230, 0.2722420, 0.7630580, 0.2540140, 0.3949320, 0.8749370, 0.7969770, 0.5023590, 0.1011950, 0.7927850, 0.4276220, 0.5525170, 0.4009600, 0.7525120, 0.1134650, 0.1582330, 0.1724210, 0.6580450, 0.1536670, 0.3099110, 0.5972860, 0.8417020, 0.5390270, 0.9634150, 0.1598230, 0.5173500, 0.7778150, 0.0027191, 0.3903830, 0.3340860, 0.8659850, 0.8017120, 0.3431660, 0.0411105, 0.7254650, 0.6544150, 0.1989220, 0.6085040, 0.6017340, 0.5015410, 0.4659320, 0.2536780, 0.0646381, 0.5337730, 0.1835320, 0.9469850, 0.9393080, 0.9110070, 0.7955400, 0.9025810, 0.8319450, 0.7804620, 0.3488540, 0.7372440, 0.7156640, 0.2623570, 0.2192500, 0.5086040, 0.3196460, 0.2439410, 0.4706060, 0.5005380, 0.4101190, 0.1385380, 0.1257460, 0.7131290, 0.9115600, 0.2647160, 0.3115150, 0.7093650, 0.5151790, 0.1900120, 0.3008730, 0.4337210, 0.2578860, 0.7560940, 0.7533320, 0.1596150, 0.4211310, 0.9796440, 0.2532840, 0.1538850, 0.2379380, 0.8517020, 0.1628650, 0.3689910, 0.7216730, 0.2774290, 0.6483490, 0.3603420, 0.5447510, 0.1214110, 0.8483590, 0.6275330, 0.1888830, 0.6797870, 0.2426770, 0.3883020, 0.1892050, 0.6877150, 0.5114970, 0.8394800, 0.7585840, 0.3874090, 0.5029050, 0.9273580, 0.4751410, 0.0101952, 0.3012100, 0.6110530, 0.0535977, 0.5314960, 0.2409410, 0.2144790, 0.1026990, 0.8493470, 0.6862500, 0.0513688, 0.2881950, 0.9313470, 0.9163060, 0.4817980, 0.9682590, 0.3976360, 0.0303608, 0.4123950, 0.8060110, 0.6185870, 0.6782290, 0.2884480, 0.7394100, 0.9973570, 0.4181960, 0.8132300, 0.0953438, 0.8039220, 0.6261710, 0.6892290, 0.8510310, 0.8049950, 0.5868210, 0.9191750, 0.5229240, 0.6640720, 0.3804460, 0.1474500, 0.1785750, 0.9955730, 0.7466310, 0.8577100, 0.1542650, 0.3396370, 0.7599620, 0.6970790, 0.2751530, 0.3698680, 0.4625630, 0.0667386, 0.1671940, 0.9043440, 0.2553890, 0.2272860, 0.7671100, 0.6262330, 0.1687030, 0.5139800, 0.1534110, 0.2727000, 0.3386930, 0.7833380, 0.3852220, 0.3599640, 0.1193900, 0.6366530, 0.0118656, 0.6782470, 0.7041950, 0.3664410, 0.6935960, 0.7774520, 0.9623710, 0.3474920, 0.5529210, 0.1853470, 0.6368900, 0.8758950, 0.2782150, 0.8270340, 0.7486750, 0.8229390, 0.0615322, 0.7431030, 0.1281490, 0.4662780, 0.0476892, 0.8186380, 0.3395020, 0.7366790, 0.6002210, 0.6658090, 0.8097920, 0.8506350, 0.2999700, 0.7706250, 0.4492020, 0.4098420, 0.4686980, 0.3031500, 0.9270150, 0.5890420, 0.5812820, 0.1643930, 0.8799180, 0.8546590, 0.3992060, 0.3231450, 0.1411380, 0.9934300, 0.7118510, 0.6305330, 0.0196712, 0.0838786, 0.6634340, 0.5875180, 0.4966150, 0.5372050, 0.5765520, 0.9392130, 0.0729185, 0.3872140, 0.2465970, 0.2561480, 0.4646000, 0.2744950, 0.7690030, 0.5526430, 0.3487990, 0.7636040, 0.7527870, 0.6296000, 0.1216730, 0.6340800, 0.0570104, 0.1132320, 0.5980700, 0.8497360, 0.6013900, 0.2326680, 0.4597970, 0.9609830, 0.5664260, 0.7010390, 0.0587407, 0.8614670, 0.6858380, 0.4757830, 0.3554550, 0.9218950, 0.1657250, 0.1000910, 0.3528310, 0.1644170, 0.7258430, 0.1717560, 0.2065620, 0.9503600, 0.3068870, 0.1448100, 0.6543000, 0.4351800, 0.0563767, 0.5389510, 0.9185840, 0.9492810, 0.4464240, 0.0063676, 0.6555070, 0.3915380, 0.4150430, 0.7040400, 0.2247390, 0.0916648, 0.2896940, 0.7560080, 0.5595030, 0.1645240, 0.0375536, 0.3017080, 0.3744600, 0.3634720, 0.2158470, 0.2267270, 0.9446030, 0.1805900, 0.8105720, 0.9635490, 0.4157950, 0.1066380, 0.9775340, 0.3421560, 0.8292740, 0.2884450, 0.3554690, 0.1792120, 0.9298060, 0.0517262, 0.6277160, 0.5480770, 0.0270531, 0.0105302, 0.3204780, 0.7312290, 0.7706980, 0.0077944, 0.6330730, 0.8115800, 0.3443620, 0.6069900, 0.0321039, 0.2415050, 0.2931840, 0.5024290, 0.5844580, 0.8618330, 0.1763640, 0.0403794, 0.4636390, 0.9983470, 0.1433290, 0.2505820, 0.1612750, 0.6114430, 0.8235630, 0.4503700, 0.4577530, 0.3641000, 0.2849600, 0.2054730, 0.6688810, 0.1574880, 0.8190680, 0.0842486, 0.5118840, 0.0442898, 0.0719923, 0.3096410, 0.2333130, 0.4310580, 0.0744885, 0.8803740, 0.2651210, 0.6087750, 0.1337880, 0.2772760, 0.7187650, 0.8499810, 0.9713510, 0.7428380, 0.9753850, 0.4540920, 0.5991570, 0.1257440, 0.7038800, 0.9330650, 0.1176710, 0.4304660, 0.0217931, 0.5095570, 0.4615570, 0.4820450, 0.4882320, 0.4713280, 0.1966680, 0.4232040, 0.9114160, 0.3048440, 0.1762120, 0.8979470, 0.2395600, 0.4472710, 0.5340150, 0.9507420, 0.7082640, 0.3091170, 0.1599090, 0.6285780, 0.8505460, 0.6334720, 0.1088460, 0.7681180, 0.7428290, 0.3480070, 0.2275180, 0.4374250, 0.9336200, 0.8848590, 0.3796180, 0.9846750, 0.7181720, 0.3346840, 0.8877670, 0.4791620, 0.6343160, 0.4135160, 0.1445380, 0.3517390, 0.6833030, 0.1894860, 0.6559010, 0.5416060, 0.9455980, 0.0630410, 0.7894870, 0.1063730, 0.7834430, 0.5968300, 0.2194690, 0.2356460, 0.6512020, 0.1082280, 0.1583040, 0.9294810, 0.9096720, 0.2072550, 0.9272000, 0.2124000, 0.2113970, 0.1190190, 0.3542760, 0.9866460, 0.4867160, 0.4520720, 0.9646480, 0.1915560, 0.1913760, 0.1774130, 0.0905867, 0.5412160, 0.5141390, 0.3312230, 0.3897770, 0.7886660, 0.9918440, 0.1793840, 0.8219620, 0.9140640, 0.2473600, 0.7422730, 0.0175527, 0.4575920, 0.1967830, 0.2141540, 0.6821420, 0.1306720, 0.4774150, 0.9150480, 0.2154790, 0.0811664, 0.1467360, 0.1699280, 0.1883030, 0.4053590, 0.9198770, 0.3591720, 0.4220780, 0.5275850, 0.1223400, 0.6000330, 0.1642760, 0.9152380, 0.5301780, 0.0597655, 0.5298160, 0.7529510, 0.8689010, 0.9663090, 0.9860990, 0.1309810, 0.4784300, 0.3897920, 0.0165162, 0.8915030, 0.5746520, 0.3505860, 0.0048667, 0.0337861, 0.0161844, 0.5863440, 0.0721362, 0.7393140, 0.6585870, 0.3980190, 0.1139030, 0.8071320, 0.2369480, 0.1519770, 0.2686370, 0.4984640, 0.7120270, 0.7910320, 0.4800250, 0.8673780, 0.7896640, 0.4557070, 0.9781970, 0.4146930, 0.2605860, 0.6596100, 0.3621220, 0.7367160, 0.7356970, 0.5906050, 0.7040340, 0.2799910, 0.8196960, 0.8011910, 0.0933821, 0.1316560, 0.4683520, 0.1225180, 0.7037110, 0.7645390, 0.3998230, 0.0400991, 0.3153030, 0.7980700, 0.3127620, 0.4664840, 0.5857620, 0.0579393, 0.4819720, 0.8379730, 0.6985410, 0.5487800, 0.3785740, 0.4979750, 0.1178110, 0.4286530, 0.0224960, 0.6469370, 0.6678220, 0.2389980, 0.7627590, 0.4923820, 0.0902086, 0.5174950, 0.0110347, 0.4467340, 0.3727500, 0.5871650, 0.9154050, 0.7665720, 0.8959990, 0.5777870, 0.4324170, 0.3537040, 0.5121720, 0.1032680, 0.7705380, 0.3102530, 0.7680280, 0.6868090, 0.0377845, 0.2272750, 0.6938420, 0.9929090, 0.1016760, 0.7446470, 0.3260430, 0.1150130, 0.2172980, 0.1410080, 0.5312020, 0.2794450, 0.9427950, 0.0387187, 0.8092000, 0.4621480, 0.2400470, 0.8404690, 0.6400280, 0.9373180, 0.9450510, 0.1536550, 0.9085070, 0.6399940, 0.0796639, 0.3908080, 0.5089620, 0.5659390, 0.2324310, 0.1345850, 0.7597180, 0.4760650, 0.4775130, 0.8250780, 0.5362740, 0.6660880, 0.4673590, 0.1167550, 0.1183440, 0.4013680, 0.0737290, 0.6180250, 0.8281620, 0.6251810, 0.4811640, 0.8816040, 0.6076840, 0.6028220, 0.2359810, 0.0511874, 0.3943580, 0.0256890, 0.5908450, 0.2962270, 0.5649830, 0.0970786, 0.7535320, 0.5981730, 0.3255790, 0.9093880, 0.0038028, 0.1154520, 0.2973620, 0.4258280, 0.9695050, 0.1135230, 0.1592360, 0.3249330, 0.6658700, 0.3911600, 0.5663430, 0.7563530, 0.5924910, 0.0190206, 0.5038270, 0.1763310, 0.8701610, 0.8796530, 0.2447070, 0.0157126, 0.9815030, 0.3120840, 0.7245960, 0.6498620, 0.4466870, 0.2021680, 0.7144230, 0.1907990, 0.7360930, 0.8915180, 0.2733100, 0.0439463, 0.3169390, 0.0288732, 0.1470670, 0.6404400, 0.8466210, 0.3346020, 0.6630830, 0.9504630, 0.9652370, 0.1721440, 0.2331500, 0.6952910, 0.6815980, 0.1046910, 0.8366110, 0.5040770, 0.9193130, 0.3579040, 0.9858360, 0.2729790, 0.7858510, 0.2591820, 0.1081410, 0.4174980, 0.1217800, 0.1940420, 0.7993890, 0.8563220, 0.4843270, 0.7441990, 0.1465730, 0.0162954, 0.8985030, 0.2766020, 0.5578080, 0.2670190, 0.0502883, 0.2940920, 0.6173670, 0.4159100, 0.5907810, 0.2001890, 0.2175100, 0.1889170, 0.5266910, 0.4359080, 0.1240500, 0.7156460, 0.5169750, 0.5325540, 0.1932510, 0.7486910, 0.7304160, 0.6319170, 0.8614480, 0.3801180, 0.9685100, 0.1092060, 0.8712240, 0.3518500, 0.0237457, 0.7491750, 0.4444270, 0.0765558, 0.3303360, 0.7903140, 0.6653800, 0.6461970, 0.2742680, 0.6865190, 0.3039870, 0.1620540, 0.6462330, 0.0311463, 0.6533520, 0.7238770, 0.0531298, 0.8442920, 0.5958600, 0.1626840, 0.0330969, 0.4215890, 0.3691840, 0.0603153, 0.2907140, 0.3296850, 0.0680191, 0.3615490, 0.9116310, 0.5784430, 0.5083830, 0.4337940, 0.2286420, 0.8150150, 0.5595470, 0.1232180, 0.8067230, 0.3951520, 0.2058890, 0.2386480, 0.9393790, 0.1260620, 0.3820600, 0.7649190, 0.9305270, 0.4580090, 0.0003186, 0.0211318, 0.8776000, 0.9885220, 0.9450760, 0.9502250, 0.5350880, 0.9972050, 0.5984590, 0.0261845, 0.9399730, 0.3124570, 0.0272654, 0.5073800, 0.1164280, 0.8691750, 0.9911930, 0.0655040, 0.0997293, 0.8841480, 0.5807630, 0.0396459, 0.0428236, 0.7684770, 0.2667640, 0.8719890, 0.2475310, 0.1402070, 0.6717210, 0.3903170, 0.0391283, 0.5223620, 0.2058450, 0.4207270, 0.8952940, 0.6086110, 0.8657250, 0.5699930, 0.5088970, 0.8218170, 0.2570150, 0.6481870, 0.4293310, 0.2168180, 0.7483350, 0.3125680, 0.1482570, 0.6894850, 0.1114780, 0.1780420, 0.3732060, 0.4103630, 0.9342830, 0.6088270, 0.4323250, 0.1119860, 0.9970970, 0.6001310, 0.4379450, 0.6046880, 0.5495140, 0.5889430, 0.7489020, 0.0863242, 0.7324320, 0.3897080, 0.6670990, 0.3906590, 0.2663960, 0.7710760, 0.5196320, 0.5872270, 0.3432720, 0.3468280, 0.7511010, 0.3182160, 0.6993060, 0.7924660, 0.3337240, 0.4226380, 0.7607750, 0.6390950, 0.3487690, 0.6130960, 0.3756050, 0.4485050, 0.0730609, 0.4770330, 0.5642550, 0.8758830, 0.8470520, 0.3893150, 0.7947640, 0.0633266, 0.8334670, 0.7399960, 0.0903747, 0.0607952, 0.6310530, 0.3245470, 0.0370114, 0.9295440, 0.8126360, 0.5692620, 0.3452000, 0.8201940, 0.8052670, 0.7467440, 0.5630620, 0.0213251, 0.4271030, 0.3726190, 0.4939020, 0.7422050, 0.5067460, 0.8529400, 0.3609770, 0.5047280, 0.8543610, 0.7068410, 0.8400340, 0.3673990, 0.0666171, 0.1525530, 0.1853470, 0.9967570, 0.6754510, 0.6143850, 0.5820490, 0.7457650, 0.4172310, 0.1659790, 0.9973370, 0.4620050, 0.2868410, 0.2246220, 0.0639499, 0.2915940, 0.5355490, 0.4957550, 0.1985910, 0.3229670, 0.8415400, 0.1576850, 0.7456210, 0.2267380, 0.7115610, 0.8032390, 0.6952510, 0.7284160, 0.7828590, 0.1403680, 0.0417813, 0.9040710, 0.4298260, 0.6901370, 0.4318890, 0.3461010, 0.1638690, 0.4809220, 0.0433490, 0.6662620, 0.1730030, 0.9458290, 0.3255460, 0.9539980, 0.2170530, 0.3336770, 0.9894470, 0.8922120, 0.6389090, 0.1351250, 0.4352270, 0.4406590, 0.6074520, 0.7203950, 0.5575430, 0.0231393, 0.4929200, 0.9771930, 0.5234610, 0.3305440, 0.6294730, 0.1801440, 0.2433040, 0.1597350, 0.4279930, 0.6119740, 0.3598140, 0.7952550, 0.0362311, 0.3467350, 0.0273461, 0.3042900, 0.9981560, 0.1479820, 0.0337134, 0.3004260, 0.1872150, 0.5620620, 0.1467140, 0.7442870, 0.7450060, 0.2847000, 0.3859220, 0.8953330, 0.7903200, 0.4610900, 0.1110170, 0.3040630, 0.2855620, 0.6092670, 0.8389160, 0.3143070, 0.6930530, 0.3072500, 0.2487770, 0.4081040, 0.0585860, 0.3219540, 0.3871980, 0.3789600, 0.2786490, 0.3840250, 0.7661320, 0.3600480, 0.4171690, 0.7685190, 0.9781080, 0.1785640, 0.8211030, 0.3835230, 0.1483930, 0.3638810, 0.4231840, 0.9087600, 0.9789650, 0.7039440, 0.4794650, 0.6024890, 0.9027490, 0.1920950, 0.9880840, 0.5651170, 0.6956230, 0.4955580, 0.9770970, 0.0490451, 0.2778970, 0.2829820, 0.9521600, 0.6234470, 0.1411300, 0.9559110, 0.8800280, 0.6016250, 0.6803420, 0.8007560, 0.6881750, 0.7201090, 0.2476530, 0.1467040, 0.5571980, 0.0860618, 0.5251660, 0.6666060, 0.0146429, 0.5121510, 0.1989260, 0.6929840, 0.5136340, 0.2663840, 0.8539490, 0.4110460, 0.5079280, 0.6994980, 0.6839610, 0.6962420, 0.8817040, 0.6863400, 0.6569070, 0.9153400, 0.5722140, 0.9999280, 0.3001000, 0.6944590, 0.4174250, 0.0069966, 0.9186340, 0.9032210, 0.6254260, 0.3574980, 0.0139199, 0.5840910, 0.0930363, 0.0053798, 0.6759190, 0.6690280, 0.2179800, 0.7357860, 0.3412730, 0.6290360, 0.5444670, 0.0765703, 0.4649790, 0.6025890, 0.3708240, 0.0112323, 0.0511709, 0.8500810, 0.0479759, 0.8666020, 0.3800670, 0.4580730, 0.1807690, 0.3795010, 0.4794500, 0.6118290, 0.2418970, 0.4298510, 0.2177560, 0.9706920, 0.7887880, 0.8673600, 0.5141430, 0.4800150, 0.7291270, 0.3681920, 0.6654340, 0.7415560, 0.1264070, 0.2363650, 0.8725310, 0.2824560, 0.7926670, 0.1605100, 0.0208207, 0.2149490, 0.5766840, 0.2995220, 0.8751850, 0.9653430, 0.8202210, 0.8933690, 0.7001970, 0.6324680, 0.2069050, 0.4867670, 0.1235510, 0.4856790, 0.4989490, 0.6239880, 0.3966060, 0.6814500, 0.3262560, 0.1835250, 0.0673006, 0.2535210, 0.8595840, 0.4089660, 0.5532730, 0.8873600, 0.9807090, 0.0427780, 0.2486150, 0.2255140, 0.7914800, 0.7541420, 0.0677359, 0.3355470, 0.0058455, 0.5135960, 0.0050992, 0.6439750, 0.4064040, 0.6406990, 0.0142548, 0.9378280, 0.8887350, 0.7639010, 0.9711190, 0.9547240, 0.5039120, 0.1434460, 0.5478370, 0.5018390, 0.7144760, 0.4444180, 0.1657780, 0.2194200, 0.0272047, 0.5823320, 0.3275310, 0.7779070, 0.1731240, 0.0786923, 0.9885610, 0.9331250, 0.9326090, 0.0126710, 0.8182930, 0.3977710, 0.0172242, 0.0790679, 0.3038380, 0.3164670, 0.3399450, 0.8781690, 0.4689860, 0.3060240, 0.0056492, 0.5896970, 0.0854484, 0.9534870, 0.3512450, 0.4689500, 0.9404640, 0.8529460, 0.3589750, 0.8805410, 0.2612130, 0.1134680, 0.9620650, 0.9008180, 0.6519580, 0.4279030, 0.3258300, 0.7049190, 0.0530086, 0.8184050, 0.7095850, 0.4871820, 0.1760130, 0.7305800, 0.1877590, 0.2358550, 0.6174560, 0.7325930, 0.3414740, 0.9410190, 0.3203310, 0.1870220, 0.5819880, 0.1944680, 0.1162880, 0.2202780, 0.4172320, 0.9069970, 0.0983290, 0.9594200, 0.3531670, 0.8994970, 0.9516290, 0.6024680, 0.6491690, 0.1330760, 0.4079180, 0.5849880, 0.1203810, 0.3420610, 0.7381950, 0.3958660, 0.4342030, 0.1063790, 0.0718363, 0.1014690, 0.7255560, 0.3019210, 0.4826340, 0.8896090, 0.7147060, 0.6606950, 0.0331155, 0.3916920, 0.1897560, 0.2463040, 0.9364730, 0.6711940, 0.6038450, 0.1977650, 0.5897340, 0.1895180, 0.6472920, 0.9089240, 0.4307910, 0.7584440, 0.1886510, 0.2403110, 0.6542060, 0.1270170, 0.7894010, 0.2023400, 0.5314730, 0.4221230, 0.5304350, 0.5549740, 0.8045940, 0.7054910, 0.6420870, 0.7455960, 0.6143490, 0.3105300, 0.7770070, 0.6138510, 0.6947270, 0.3015500, 0.8415390, 0.6324010, 0.3603590, 0.9484740, 0.1967150, 0.2290850, 0.1385560, 0.8713360, 0.4297970, 0.7486860, 0.8457380, 0.7040300, 0.6947830, 0.9969930, 0.6491710, 0.5692650, 0.9386200, 0.7367540, 0.5729650, 0.6603930, 0.5096410, 0.1811190, 0.0607770, 0.8775210, 0.0572442, 0.0776710, 0.3638410, 0.8144830, 0.2982850, 0.3827090, 0.0757509, 0.2552840, 0.7774080, 0.1171280, 0.2684520, 0.0155161, 0.3328260, 0.5197210, 0.1690260, 0.2943240, 0.5541910, 0.6372290, 0.1800880, 0.8936980, 0.0180155, 0.2527280, 0.9077520, 0.4667450, 0.8383220, 0.0487360, 0.0310284, 0.9932800, 0.6723090, 0.9284490, 0.1678230, 0.5622060, 0.0893037, 0.2117600, 0.4152690, 0.6480720, 0.0392260, 0.1355680, 0.5672940, 0.7648580, 0.0244483, 0.5497980, 0.6115290, 0.7835850, 0.3296290, 0.8402310, 0.0909212, 0.1196230, 0.2172090, 0.0367870, 0.0201069, 0.8331920, 0.3046530, 0.5010090, 0.3373540, 0.5362650, 0.0484083, 0.4592430, 0.1711040, 0.3684340, 0.0674122, 0.6697130, 0.5678630, 0.2765720, 0.0428114, 0.9859250, 0.7011220, 0.4544730, 0.9023530, 0.9650260, 0.6050220, 0.4184570, 0.8243910, 0.5423950, 0.6709940, 0.7867750, 0.3756660, 0.8181140, 0.7518750, 0.2384630, 0.9127780, 0.3950750, 0.1901880, 0.9306440, 0.2685280, 0.3881180, 0.4799110, 0.1028810, 0.3955570, 0.5580840, 0.4043070, 0.7344720, 0.8851670, 0.7386420, 0.9016370, 0.0648124, 0.2893720, 0.9755750, 0.1575880, 0.6717530, 0.9305470, 0.6787240, 0.7284680, 0.1059990, 0.4720460, 0.8299130, 0.8837900, 0.3565200, 0.2417760, 0.9895820, 0.6927380, 0.9032660, 0.3966060, 0.4380030, 0.6052570, 0.3503200, 0.4241050, 0.0996658, 0.3851940, 0.7718420, 0.2052060, 0.6069690, 0.5070080, 0.9241850, 0.5953750, 0.7103970, 0.8788110, 0.9603380, 0.9950640, 0.6578640, 0.2818210, 0.2792460, 0.1440100, 0.3124180, 0.5928510, 0.6361660, 0.5018210, 0.5920670, 0.2476340, 0.1881220, 0.2462910, 0.6007210, 0.7450060, 0.2713220, 0.7658820, 0.0786912, 0.4894550, 0.3971030, 0.1232920, 0.1844170, 0.6630790, 0.2277350, 0.1555700, 0.2906220, 0.3708960, 0.7748850, 0.4161810, 0.9736690, 0.1509800, 0.2140620, 0.8982070, 0.4415930, 0.1494230, 0.1604290, 0.1990320, 0.1556970, 0.6089220, 0.4599240, 0.1748290, 0.9641130, 0.0709676, 0.8187310, 0.8006890, 0.0961359, 0.9981690, 0.4695020, 0.9861410, 0.8710280, 0.1079930, 0.5411980, 0.0856880, 0.1831780, 0.5552190, 0.2614090, 0.9925410, 0.6715800, 0.0767847, 0.7883510, 0.9304150, 0.3383720, 0.2465090, 0.8398170, 0.3750660, 0.0895940, 0.1413190, 0.3773660, 0.4449410, 0.2547200, 0.7371920, 0.7530190, 0.3361020, 0.8517140, 0.5220190, 0.3963820, 0.8799920, 0.8306800, 0.7261260, 0.9946910, 0.2147760, 0.7709730, 0.8286000, 0.0657721, 0.4232100, 0.0323970, 0.5957580, 0.2198150, 0.2475880, 0.0903869, 0.9304430, 0.8871300, 0.7907850, 0.1501000, 0.6285370, 0.0060634, 0.7585790, 0.8413310, 0.7645360, 0.0822761, 0.7858810, 0.3962700, 0.8370230, 0.6224120, 0.0345241, 0.4738160, 0.9651350, 0.8012460, 0.9131650, 0.0191692, 0.9711820, 0.0219913, 0.0951320, 0.8413700, 0.3836820, 0.4464120, 0.0004582, 0.2216450, 0.6371200, 0.5107580, 0.1032810, 0.7234490, 0.4112400, 0.4562670, 0.7025890, 0.8904710, 0.1731600, 0.3472820, 0.0360796, 0.1476720, 0.6466280, 0.7381020, 0.9162220, 0.7401260, 0.0706535, 0.1229500, 0.0816709, 0.0385719, 0.9418780, 0.8254270, 0.1612520, 0.6694980, 0.5326700, 0.3422820, 0.8843840, 0.1859500, 0.3471280, 0.8734000, 0.6224260, 0.4951510, 0.9967480, 0.9686550, 0.8980860, 0.4112470, 0.0017922, 0.2290070, 0.1694690, 0.4733220, 0.0407952, 0.5809990, 0.6133650, 0.3009510, 0.3598410, 0.1003260, 0.5952380, 0.6329630, 0.5825250, 0.8062360, 0.8533290, 0.0609160, 0.4587170, 0.5693570, 0.8477520, 0.3367180, 0.7857680, 0.6896250, 0.4158170, 0.3430210, 0.6596920, 0.4187860, 0.4709480, 0.1333390, 0.1516480, 0.3537290, 0.7980220, 0.1081500, 0.8836680, 0.6461660, 0.5223790, 0.2761070, 0.0799563, 0.1726850, 0.6235330, 0.4053230, 0.4382230, 0.7259790, 0.6841380, 0.9491600, 0.9440170, 0.3841210, 0.2012550, 0.2181970, 0.2525320, 0.5962360, 0.8177800, 0.2232980, 0.2125470, 0.8238980, 0.6599280, 0.4566500, 0.7460410, 0.5067340, 0.9887100, 0.6864220, 0.3653500, 0.2436660, 0.3589200, 0.4512840, 0.0981289, 0.9952630, 0.7236670, 0.7218310, 0.8099730, 0.8141110, 0.9887400, 0.3922100, 0.3410160, 0.6213950, 0.3192930, 0.0964344, 0.6780420, 0.6123280, 0.3960160, 0.2985460, 0.5157480, 0.9437350, 0.9951450, 0.5716220, 0.1468700, 0.2902680, 0.0100090, 0.5867380, 0.0584274, 0.8069500, 0.1865340, 0.0137096, 0.8052840, 0.4502750, 0.6568890, 0.8587270, 0.2825100, 0.5080080, 0.5363220, 0.9379320, 0.2353310, 0.3441460, 0.9997060, 0.6225000, 0.0001136, 0.2379860, 0.0933501, 0.9466700, 0.5149690, 0.4348670, 0.8388820, 0.4981010, 0.0544689, 0.1428880, 0.9956100, 0.7031210, 0.1120100, 0.5791090, 0.6189760, 0.4995210, 0.8266950, 0.9720830, 0.3735180, 0.4054890, 0.1895980, 0.6411080, 0.3513720, 0.8349690, 0.9464330, 0.8212030, 0.7119760, 0.0347150, 0.6927050, 0.7287130, 0.9279290, 0.0423214, 0.5419080, 0.0986794, 0.4395800, 0.6631510, 0.3785480, 0.3959410, 0.0700278, 0.6860040, 0.2179950, 0.8194610, 0.4541530, 0.3804900, 0.3469490, 0.2169750, 0.7338240, 0.4782950, 0.4095440, 0.2806940, 0.6422090, 0.3591400, 0.6295210, 0.6837450, 0.7622400, 0.2969340, 0.6747920, 0.1082900, 0.5555310, 0.0449378, 0.2434720, 0.1776680, 0.1655840, 0.9875580, 0.4924570, 0.5931880, 0.6007370, 0.6213000, 0.9206760, 0.0385422, 0.9967580, 0.3842650, 0.4535770, 0.4689990, 0.3895050, 0.2753740, 0.4716120, 0.5136250, 0.2250340, 0.9581980, 0.5415070, 0.3758220, 0.5395650, 0.9436090, 0.4718200, 0.2130470, 0.6446440, 0.9376610, 0.8396630, 0.2134240, 0.0436052, 0.5881990, 0.6874030, 0.6994340, 0.0650040, 0.5948690, 0.6979020, 0.8709610, 0.7062200, 0.5259550, 0.5782950, 0.5778630, 0.9430990, 0.7090380, 0.1764230, 0.8807730, 0.7788570, 0.1912720, 0.6618190, 0.3337820, 0.1376100, 0.6570980, 0.3491980, 0.6732240, 0.6157340, 0.1420850, 0.5665280, 0.1392500, 0.2900810, 0.4995430, 0.6348700, 0.3859260, 0.8427740, 0.3056520, 0.8501110, 0.4894240, 0.9867720, 0.0467864, 0.7659000, 0.3732920, 0.8248970, 0.0232419, 0.7279180, 0.0514450, 0.4195700, 0.5388530, 0.2600290, 0.0062874, 0.6006990, 0.7447220, 0.8328340, 0.8330300, 0.0622784, 0.1231960, 0.1390060, 0.9285450, 0.6658350, 0.0013372, 0.8372210, 0.2017380, 0.4500200, 0.5746080, 0.1850240, 0.6078430, 0.6243930, 0.8957720, 0.3742210, 0.3851430, 0.6317150, 0.9887470, 0.6447660, 0.8945110, 0.6217990, 0.1178140, 0.7991900, 0.9277560, 0.2355290, 0.5509700, 0.8306270, 0.7471910, 0.7010700, 0.9324260, 0.5962370, 0.0918996, 0.1852300, 0.8266290, 0.5952830, 0.2989090, 0.7255950, 0.8108870, 0.6781480, 0.5605800, 0.8817860, 0.9128430, 0.6225460, 0.0373080, 0.6764460, 0.2307220, 0.2484460, 0.5394630, 0.7784840, 0.4441150, 0.2333820, 0.4341850, 0.5277350, 0.8043690, 0.4155310, 0.4089220, 0.5546250, 0.7866070, 0.0593978, 0.2544930, 0.8899290, 0.2612840, 0.1087990, 0.6243820, 0.2405500, 0.5056270, 0.8609370, 0.7865130, 0.7699840, 0.6513300, 0.7076120, 0.8798100, 0.4117680, 0.5533810, 0.7277270, 0.3234570, 0.2296480, 0.1483080, 0.9620880, 0.9870980, 0.2134340, 0.8936250, 0.4997170, 0.3966200, 0.3905010, 0.0779684, 0.3100650, 0.2004820, 0.6716580, 0.1090680, 0.7277720, 0.9077130, 0.3031230, 0.7938920, 0.6619360, 0.9126580, 0.2993680, 0.0976682, 0.2096540, 0.3557550, 0.6906320, 0.0192524, 0.8001940, 0.9493270, 0.6600840, 0.3180520, 0.2776060, 0.0456789, 0.1643590, 0.1263820, 0.4981630, 0.5531860, 0.6460530, 0.9153240, 0.3262450, 0.9060420, 0.4381480, 0.2655070, 0.6220110, 0.7731080, 0.0746926, 0.3258660, 0.6195530, 0.0238042, 0.0494728, 0.5469910, 0.6486250, 0.2046000, 0.1811620, 0.7433750, 0.1971430, 0.9528520, 0.0372530, 0.9945320, 0.0483653, 0.1318760, 0.1382750, 0.4316350, 0.6735530, 0.5703900, 0.5071450, 0.5146910, 0.9566450, 0.7993770, 0.0072045, 0.2289590, 0.4828670, 0.4713780, 0.6267050, 0.9567290, 0.5322800, 0.3992350, 0.0414665, 0.2177130, 0.0675323, 0.4371870, 0.6389060, 0.9117010, 0.4611630, 0.4987740, 0.9435350, 0.7917080, 0.2329080, 0.8987710, 0.0662942, 0.9859900, 0.9286290, 0.0784090, 0.4422350, 0.5743120, 0.5492650, 0.0503034, 0.2426240, 0.4299090, 0.0313762, 0.7736040, 0.7539990, 0.6163010, 0.9190020, 0.7617990, 0.1596090, 0.4195720, 0.3428710, 0.1537420, 0.4025830, 0.5549030, 0.1794270, 0.9804720, 0.2876570, 0.8771020, 0.9514760, 0.9566950, 0.7846510, 0.5104040, 0.4382130, 0.9296160, 0.5140710, 0.3999790, 0.3547810, 0.7662460, 0.1970510, 0.0823942, 0.2023180, 0.0875088, 0.7351980, 0.0461193, 0.5386040, 0.1650630, 0.5871850, 0.0838942, 0.5754930, 0.1493490, 0.8660350, 0.4174760, 0.5550900, 0.2649170, 0.9829610, 0.9645240, 0.4089480, 0.4492080, 0.9485910, 0.6514310, 0.8420370, 0.6669190, 0.2831850, 0.6100210, 0.6843430, 0.9210000, 0.9360520, 0.4253090, 0.7688450, 0.2573410, 0.3576130, 0.6624220, 0.0223378, 0.4504170, 0.8579240, 0.5716350, 0.8877150, 0.6968320, 0.6980030, 0.4596540, 0.5645860, 0.5228780, 0.1846030, 0.4036370, 0.1589910, 0.3562170, 0.6240300, 0.8243120, 0.6425490, 0.6881200, 0.5492300, 0.2165940, 0.4401810, 0.2937890, 0.1139720, 0.0617991, 0.8881820, 0.2263540, 0.9391910, 0.7108330, 0.8636930, 0.1801000, 0.9987580, 0.8577810, 0.6482310, 0.7912210, 0.2120850, 0.9524890, 0.4876490, 0.0689676, 0.4478100, 0.1701700, 0.9575700, 0.5005050, 0.4650070, 0.2746510, 0.5426360, 0.2314290, 0.7362720, 0.8333800, 0.8473660, 0.5771190, 0.8354910, 0.6755110, 0.5796710, 0.1455490, 0.6810120, 0.2005480, 0.7653910, 0.8236300, 0.5022740, 0.4030360, 0.5002000, 0.8318800, 0.6395140, 0.7729650, 0.8780780, 0.3223330, 0.7665420, 0.6465510, 0.2142010, 0.2494030, 0.5218690, 0.5230330, 0.8718470, 0.9528840, 0.5890740, 0.5312180, 0.6196740, 0.5860810, 0.8318770, 0.9138940, 0.0869406, 0.4862420, 0.6019470, 0.4304760, 0.5695200, 0.7386110, 0.2835530, 0.2321850, 0.7336260, 0.1303520, 0.6225520, 0.4601160, 0.0719695, 0.0806398, 0.5310520, 0.0537306, 0.3360890, 0.2552100, 0.8637270, 0.4395860, 0.5413240, 0.8957090, 0.5834730, 0.5526150, 0.3347890, 0.6834370, 0.9157390, 0.0278103, 0.1773640, 0.2769210, 0.8403520, 0.0732345, 0.4421500, 0.1814370, 0.7561590, 0.0596628, 0.8754340, 0.4598350, 0.1145160, 0.5617220, 0.7965560, 0.3213860, 0.9305710, 0.5932510, 0.2554210, 0.7970890, 0.6595630, 0.5520270, 0.6741260, 0.7050550, 0.0838225, 0.9061960, 0.4797790, 0.5792300, 0.4570110, 0.8775860, 0.1758590, 0.7862640, 0.0338609, 0.7451920, 0.5468650, 0.7827510, 0.0849230, 0.1298060, 0.8379770, 0.5031850, 0.8276640, 0.6819890, 0.4249230, 0.2598000, 0.1157770, 0.6068930, 0.5740890, 0.4415440, 0.1819040, 0.2745940, 0.3181970, 0.7538600, 0.4897830, 0.7767980, 0.4303860, 0.5372660, 0.1890400, 0.9807920, 0.1804500, 0.0124766, 0.0992348, 0.9438720, 0.0056217, 0.7304820, 0.8932080, 0.6067380, 0.9939170, 0.1524180, 0.1192620, 0.9534120, 0.4624660, 0.4133580, 0.0710641, 0.2693850, 0.8794040, 0.6497530, 0.8657430, 0.5933900, 0.5652140, 0.8555440, 0.1647700, 0.4761950, 0.5948740, 0.9978250, 0.7217750, 0.0260677, 0.4716110, 0.4297860, 0.0234541, 0.3417860, 0.3559310, 0.0207681, 0.6615400, 0.1397110, 0.0843639, 0.0389179, 0.5408660, 0.0014189, 0.0482221, 0.7750620, 0.6956560, 0.0380432, 0.4552230, 0.6604860, 0.5838500, 0.1833700, 0.1961200, 0.1357790, 0.8624990, 0.5192630, 0.1524650, 0.0195962, 0.7480690, 0.3595640, 0.1296710, 0.9679720, 0.4713160, 0.1682010, 0.2227430, 0.1930720, 0.0171584, 0.0000297, 0.1169670, 0.8566750, 0.9947340, 0.2438990, 0.6417860, 0.9970170, 0.2551050, 0.3774420, 0.9567540, 0.5661170, 0.0686075, 0.7774380, 0.2294500, 0.1857090, 0.1011480, 0.2455830, 0.2845490, 0.1686530, 0.4258630, 0.0006054, 0.3003460, 0.1454000, 0.9397850, 0.5922710, 0.5993330, 0.0516510, 0.3089320, 0.8713440, 0.9055200, 0.1225540, 0.1115020, 0.1242590, 0.7533290, 0.7835850, 0.7370980, 0.9488810, 0.1990900, 0.3276610, 0.3197010, 0.8997530, 0.4672240, 0.2972340, 0.6190850, 0.3034990, 0.7573440, 0.9176880, 0.3372250, 0.9590420, 0.5254920, 0.8786890, 0.0814828, 0.8283510, 0.7414630, 0.7915840, 0.6760600, 0.7470000, 0.6184570, 0.9265100, 0.8392790, 0.9279440, 0.4855950, 0.5865210, 0.3162620, 0.4468860, 0.8674150, 0.0723330, 0.6608350, 0.7163320, 0.6446970, 0.7793210, 0.6205150, 0.2355320, 0.3098320, 0.4793850, 0.2699760, 0.1510580, 0.6900530, 0.4942870, 0.5255220, 0.2592470, 0.0920559, 0.5789040, 0.8057880, 0.1724520, 0.4202140, 0.1504980, 0.9886860, 0.9240910, 0.3300690, 0.9667350, 0.1516330, 0.2994450, 0.3425350, 0.6195060, 0.7771810, 0.2811440, 0.8740350, 0.6103830, 0.1986260, 0.6770440, 0.7772070, 0.1221080, 0.7311630, 0.9261990, 0.2640270, 0.3007460, 0.1239890, 0.1911690, 0.2403280, 0.8926990, 0.4932740, 0.8901390, 0.4293970, 0.6621970, 0.0086421, 0.7065520, 0.1144620, 0.6749230, 0.4157570, 0.5110020, 0.0733922, 0.7166840, 0.4217820, 0.2508360, 0.5285200, 0.0763232, 0.3283820, 0.4553310, 0.8396110, 0.9867340, 0.6702810, 0.0793354, 0.5027880, 0.6093780, 0.5602800, 0.0385776, 0.7720790, 0.5968190, 0.8510350, 0.4834750, 0.9949090, 0.3349500, 0.5527920, 0.1515080, 0.9158020, 0.0314329, 0.1472120, 0.0306481, 0.5613660, 0.7807330, 0.8267480, 0.4511830, 0.0210884, 0.4693850, 0.5123700, 0.3561350, 0.0155336, 0.3102680, 0.0462573, 0.5588050, 0.6182400, 0.8312270, 0.6806390, 0.0649116, 0.4419850, 0.4020650, 0.6752150, 0.4898630, 0.1998020, 0.5218660, 0.6955040, 0.2344600, 0.3694830, 0.9268360, 0.7396140, 0.4139640, 0.6611340, 0.0704857, 0.1668530, 0.2188590, 0.3637190, 0.4092210, 0.0993976, 0.5616250, 0.2968460, 0.3213100, 0.9594280, 0.1660610, 0.0012358, 0.1064200, 0.9589600, 0.8847850, 0.4269380, 0.6893990, 0.6803830, 0.6460370, 0.8565900, 0.2050320, 0.7544980, 0.7722080, 0.9120930, 0.5760500, 0.1653240, 0.3601270, 0.6979470, 0.9134320, 0.0391862, 0.6415980, 0.7453740, 0.7562730, 0.3947930, 0.5955380, 0.3000310, 0.9786780, 0.5254850, 0.5939600, 0.2188540, 0.7615720, 0.0892903, 0.8285970, 0.8887690, 0.4875750, 0.4490600, 0.7824080, 0.2600050, 0.4287540, 0.3156330, 0.3882530, 0.0825128, 0.8337650, 0.7463260, 0.1817930, 0.6291800, 0.2926390, 0.4891860, 0.1671140, 0.0728832, 0.2652410, 0.2256680, 0.5969140, 0.5380120, 0.9669000, 0.4166900, 0.0548623, 0.7531170, 0.1289380, 0.8351970, 0.2806340, 0.4434640, 0.0349240, 0.6883790, 0.2735750, 0.7209020, 0.3233360, 0.6828770, 0.3456760, 0.0203226, 0.5947440, 0.3408130, 0.7342990, 0.6427410, 0.4127860, 0.9348570, 0.4328400, 0.2077800, 0.5879650, 0.1302060, 0.0557942, 0.4314490, 0.8609740, 0.7719660, 0.0310646, 0.3092130, 0.6310530, 0.7309780, 0.1673270, 0.1566830, 0.9325030, 0.4624620, 0.2914760, 0.3806410, 0.4054330, 0.4199090, 0.0471368, 0.9505160, 0.8973470, 0.3053270, 0.2756150, 0.8037170, 0.9458780, 0.2359990, 0.3735270, 0.3443220, 0.2000660, 0.6192990, 0.9502450, 0.1828130, 0.2964260, 0.0073840, 0.0528837, 0.1679100, 0.9057360, 0.3607820, 0.4331260, 0.3216090, 0.6785660, 0.7981000, 0.8494770, 0.1645380, 0.0955005, 0.8200300, 0.3715600, 0.4346330, 0.8469630, 0.4850210, 0.8464270, 0.4359500, 0.2287780, 0.6984460, 0.9774020, 0.2457150, 0.1047970, 0.6961860, 0.6525810, 0.7297550, 0.7690350, 0.5314160, 0.4153840, 0.3668830, 0.0452473, 0.6284660, 0.7929860, 0.9044870, 0.3426180, 0.0908378, 0.0012386, 0.0942077, 0.3759710, 0.9847310, 0.5850790, 0.9067570, 0.4669840, 0.2004450, 0.9001790, 0.5250550, 0.0284720, 0.7591180, 0.8129660, 0.8655630, 0.3567010, 0.0619191, 0.1995200, 0.5426200, 0.3890610, 0.5421080, 0.0127046, 0.5047470, 0.9547200, 0.9441040, 0.7976050, 0.0756759, 0.4340340, 0.1302350, 0.7470930, 0.3725870, 0.5887930, 0.0649110, 0.7808830, 0.4076440, 0.1167230, 0.8844310, 0.2890610, 0.0163426, 0.6029860, 0.6781140, 0.3520170, 0.3842390, 0.2324780, 0.9627240, 0.9869630, 0.3112890, 0.4278370, 0.2539240, 0.1001690, 0.4749090, 0.7749420, 0.6152920, 0.7716700, 0.9465580, 0.8580680, 0.7569610, 0.6919150, 0.2948180, 0.2270350, 0.4837290, 0.1255930, 0.1300670, 0.2159630, 0.7940260, 0.0668822, 0.3748260, 0.2920870, 0.2102270, 0.3421990, 0.9363280, 0.6946680, 0.5173280, 0.0237026, 0.7331400, 0.9794040, 0.8633340, 0.8894680, 0.9460880, 0.9708600, 0.2560290, 0.3227970, 0.1160650, 0.3478670, 0.4285350, 0.5304920, 0.4711310, 0.0074282, 0.5141130, 0.9874650, 0.3489480, 0.9225300, 0.7205660, 0.2915160, 0.5759680, 0.0779067, 0.3796440, 0.2503890, 0.2904310, 0.7632870, 0.3645170, 0.3265030, 0.3328770, 0.2598460, 0.2149570, 0.2936440, 0.0811037, 0.0987757, 0.1764970, 0.3905650, 0.9785400, 0.1055890, 0.7346560, 0.4089790, 0.8062540, 0.2038070, 0.8374330, 0.9029180, 0.4737750, 0.4980170, 0.6236230, 0.1704160, 0.9859470, 0.7516510, 0.3521450, 0.9143110, 0.8362350, 0.3418470, 0.7303780, 0.4589510, 0.3406170, 0.9718480, 0.2630650, 0.8321520, 0.8107230, 0.1366660, 0.2189270, 0.9460130, 0.6028200, 0.4521830, 0.1000690, 0.6194770, 0.4092530, 0.1597630, 0.7078520, 0.4898250, 0.7034910, 0.1214870, 0.9680830, 0.5107510, 0.5437780, 0.3122210, 0.3425360, 0.4319980, 0.2848010, 0.7637380, 0.0066204, 0.8210580, 0.8612910, 0.6084150, 0.5206000, 0.4000160, 0.2013460, 0.2089110, 0.1133130, 0.4874110, 0.0396798, 0.0298271, 0.4193550, 0.8367570, 0.8971670, 0.4590820, 0.7579430, 0.0554748, 0.8864810, 0.0655904, 0.7042930, 0.4489130, 0.6271160, 0.7257880, 0.1815520, 0.5070960, 0.1096480, 0.2159700, 0.1524390, 0.8178260, 0.6414290, 0.5487400, 0.2545620, 0.4438770, 0.4935160, 0.2868910, 0.7493700, 0.9447320, 0.8586320, 0.0381717, 0.3916870, 0.7028010, 0.9561550, 0.0610182, 0.2931190, 0.7662660, 0.2947690, 0.6170700, 0.3949300, 0.7763640, 0.3141540, 0.7039000, 0.3617010, 0.9535440, 0.4674720, 0.0610321, 0.1775190, 0.5328880, 0.2213340, 0.7313870, 0.9812160, 0.8361810, 0.8706710, 0.9793090, 0.8799270, 0.7783400, 0.3893790, 0.0096413, 0.7763840, 0.3894720, 0.9762850, 0.2500640, 0.6855370, 0.9384780, 0.3760090, 0.1212420, 0.2144110, 0.2584050, 0.8555530, 0.6430040, 0.7785000, 0.8367710, 0.8497650, 0.5756550, 0.5126930, 0.6716040, 0.2271960, 0.6530460, 0.9882950, 0.4913390, 0.0809872, 0.6629040, 0.5597960, 0.0032655, 0.5155890, 0.2158570, 0.4848780, 0.7150510, 0.1762830, 0.4040920, 0.8073570, 0.2543850, 0.5915800, 0.2410530, 0.9991790, 0.1935050, 0.9545450, 0.5525480, 0.0515840, 0.9183460, 0.2341990, 0.5383290, 0.4562880, 0.0378786, 0.1132200, 0.5677770, 0.2889770, 0.5436280, 0.0178214, 0.5821380, 0.9743550, 0.5644070, 0.8844180, 0.0752698, 0.8232570, 0.6152060, 0.9119230, 0.7925900, 0.5214170, 0.4475950, 0.8943800, 0.4832640, 0.2007860, 0.2346720, 0.6890510, 0.1299940, 0.3198810, 0.9554090, 0.5585450, 0.4748380, 0.8661450, 0.9529510, 0.1574180, 0.4949130, 0.8289870, 0.6707610, 0.9844790, 0.7495480, 0.3470180, 0.8367240, 0.1751030, 0.0883757, 0.6125620, 0.4248050, 0.2200380, 0.8551470, 0.7224970, 0.5970400, 0.4571160, 0.6561380, 0.3813030, 0.5198230, 0.9288880, 0.2798140, 0.2103820, 0.2751640, 0.5930750, 0.4504240, 0.4725440, 0.3923460, 0.1348060, 0.9159470, 0.9813540, 0.5437720, 0.4679860, 0.8415040, 0.4452630, 0.0811758, 0.5851860, 0.3647600, 0.3263120, 0.8667140, 0.8755910, 0.8276620, 0.4832920, 0.8253340, 0.1790770, 0.9810350, 0.3111270, 0.4229740, 0.5586630, 0.3574540, 0.0640596, 0.6098540, 0.6220120, 0.9297170, 0.3382790, 0.8300540, 0.1584870, 0.6277660, 0.6353010, 0.7085910, 0.5371470, 0.6483860, 0.9682170, 0.0451543, 0.3771620, 0.6603230, 0.6069500, 0.3851590, 0.8498530, 0.1329190, 0.6442820, 0.7640150, 0.6616630, 0.9055980, 0.0752273, 0.4395180, 0.4952400, 0.5490810, 0.8265080, 0.7455000, 0.0788394, 0.6265490, 0.7855420, 0.1977370, 0.5546790, 0.2237820, 0.2082940, 0.7199990, 0.3522380, 0.2161740, 0.6730220, 0.5069670, 0.6193560, 0.4039000, 0.6528800, 0.6198020, 0.8494710, 0.3936270, 0.4720020, 0.4667330, 0.8111860, 0.6613030, 0.4356850, 0.0414877, 0.1332240, 0.9304400, 0.4343010, 0.2846120, 0.0846275, 0.3327890, 0.9220170, 0.9247390, 0.1399950, 0.5717180, 0.5105430, 0.2336020, 0.5178130, 0.8552280, 0.2016260, 0.1767370, 0.0799954, 0.1768330, 0.8836920, 0.2355660, 0.7699420, 0.1964900, 0.6619890, 0.1499400, 0.8205310, 0.0902560, 0.1245180, 0.4341200, 0.7510990, 0.3467640, 0.1529500, 0.9069330, 0.2900590, 0.0751384, 0.3831170, 0.3743330, 0.0984511, 0.2463880, 0.2120980, 0.9201260, 0.2268060, 0.8718570, 0.5609560, 0.1865460, 0.4587110, 0.5859730, 0.3084270, 0.8764780, 0.4858410, 0.3677510, 0.2925180, 0.4643840, 0.1730460, 0.8909200, 0.1449090, 0.9308810, 0.6818370, 0.1851150, 0.2572850, 0.5734910, 0.3041700, 0.1753640, 0.9370110, 0.9941270, 0.4839090, 0.3843270, 0.2421740, 0.5509110, 0.3468110, 0.6976160, 0.2266280, 0.3526500, 0.0236813, 0.0568918, 0.8277600, 0.5543360, 0.9673210, 0.3050300, 0.3619880, 0.2377050, 0.6309850, 0.6638950, 0.9194260, 0.5500350, 0.6656070, 0.2054280, 0.4089360, 0.7104900, 0.4974710, 0.4361340, 0.0488055, 0.6103780, 0.6611150, 0.2875570, 0.4829110, 0.9006820, 0.1399710, 0.8240180, 0.3319710, 0.7583720, 0.7679350, 0.7189570, 0.5886420, 0.9166580, 0.9654170, 0.4508570, 0.6447500, 0.9883240, 0.1461130, 0.6281360, 0.4534260, 0.1395890, 0.7251240, 0.1703250, 0.8786950, 0.0235274, 0.4949860, 0.0291311, 0.8665560, 0.5056190, 0.1272090, 0.0539065, 0.9459060, 0.9001830, 0.2055900, 0.7201230, 0.7905130, 0.1696390, 0.1432770, 0.3817670, 0.7587030, 0.3999180, 0.3926660, 0.3384730, 0.0284238, 0.2984400, 0.8468680, 0.5765150, 0.5350010, 0.4431850, 0.1603970, 0.7269900, 0.9516220, 0.5233250, 0.1156910, 0.8638350, 0.5142250, 0.4983100, 0.6710690, 0.2001380, 0.8612880, 0.7801040, 0.7648210, 0.7621930, 0.5064220, 0.3788370, 0.7860140, 0.4843810, 0.6239260, 0.5404240, 0.0006382, 0.8129360, 0.9119700, 0.0227581, 0.7512380, 0.5387880, 0.3370540, 0.3841880, 0.1948490, 0.7249480, 0.9887960, 0.7846160, 0.6198900, 0.1224710, 0.9721160, 0.5880490, 0.7715780, 0.1368360, 0.5357280, 0.3863570, 0.1150800, 0.0556017, 0.9721820, 0.1042820, 0.7296220, 0.8318550, 0.2819750, 0.2123680, 0.7908470, 0.2487180, 0.6098440, 0.8081870, 0.4931930, 0.2245120, 0.2375400, 0.0250251, 0.0158882, 0.2770480, 0.2545420, 0.0564164, 0.7938120, 0.9609460, 0.8750850, 0.1094370, 0.6171970, 0.5197760, 0.2971520, 0.3807040, 0.6473100, 0.1093550, 0.5784530, 0.0481793, 0.8049220, 0.7507370, 0.9893150, 0.3517340, 0.8287500, 0.0412061, 0.2787000, 0.8891320, 0.3336770, 0.5148340, 0.6937780, 0.3731950, 0.1689270, 0.3456020, 0.3739970, 0.1019460, 0.7683310, 0.7008160, 0.4671910, 0.0400199, 0.2659930, 0.3057800, 0.3217990, 0.6705110, 0.2916020, 0.2127380, 0.6161670, 0.1699170, 0.1562050, 0.2345230, 0.8494070, 0.8323230, 0.9155160, 0.9443480, 0.6026500, 0.0760167, 0.1996820, 0.9554680, 0.6878040, 0.3395310, 0.0013971, 0.0761547, 0.1714670, 0.7786540, 0.4118640, 0.3731030, 0.2223350, 0.4865000, 0.6337310, 0.9400140, 0.1610940, 0.0116855, 0.9413800, 0.3768320, 0.5477960, 0.1478770, 0.6730070, 0.3834410, 0.7447030, 0.9742050, 0.8254200, 0.5398490, 0.1323470, 0.8805620, 0.7466560, 0.6467550, 0.4304130, 0.9486190, 0.1328520, 0.4668080, 0.9334420, 0.0849821, 0.2555340, 0.1704170, 0.9072950, 0.4479820, 0.2276410, 0.7551440, 0.1697240, 0.7004370, 0.2989380, 0.1194520, 0.1012210, 0.0781414, 0.8208570, 0.5873560, 0.2032170, 0.8211250, 0.6263520, 0.5511560, 0.4855460, 0.6859220, 0.3359880, 0.7101460, 0.9778610, 0.8629300, 0.4846240, 0.9019890, 0.3937970, 0.8822800, 0.9620730, 0.0864188, 0.9301350, 0.6495690, 0.2602090, 0.4641930, 0.4681950, 0.6260900, 0.9400910, 0.9155740, 0.5473920, 0.2659020, 0.1374720, 0.8277920, 0.9650370, 0.2758160, 0.8952720, 0.6121050, 0.0354861, 0.8549950, 0.8946600, 0.7142390, 0.7874850, 0.3405000, 0.8207900, 0.7906770, 0.9477660, 0.8946680, 0.1484060, 0.2379060, 0.0854444, 0.4259210, 0.2797500, 0.1692910, 0.9502210, 0.6813660, 0.2945520, 0.6172130, 0.1426570, 0.9706440, 0.6434470, 0.3346330, 0.7674170, 0.1548520, 0.2705400, 0.9523350, 0.3900370, 0.0903934, 0.1192310, 0.8141470, 0.7262670, 0.1629230, 0.1795430, 0.2611120, 0.1528900, 0.0300276, 0.6520350, 0.1756130, 0.0508901, 0.6659140, 0.5332550, 0.2521160, 0.8225930, 0.7993850, 0.5004140, 0.3307460, 0.2208050, 0.4726510, 0.4923430, 0.5026430, 0.0132745, 0.1848080, 0.1072270, 0.9110430, 0.0882753, 0.7899890, 0.3133580, 0.0426921, 0.6841230, 0.5331850, 0.7254690, 0.8913450, 0.9923520, 0.6926320, 0.6678360, 0.8451710, 0.5333120, 0.6991220, 0.0577702, 0.3836210, 0.9620800, 0.1023540, 0.7088660, 0.9802860, 0.2026860, 0.8280000, 0.3479380, 0.2375370, 0.2170530, 0.2327360, 0.5243760, 0.3814580, 0.4173100, 0.8747960, 0.9721930, 0.0236887, 0.1815610, 0.4373740, 0.4203510, 0.5702380, 0.9979320, 0.6528210, 0.7459620, 0.9332860, 0.0866012, 0.9670140, 0.5707320, 0.3524230, 0.0321593, 0.7395670, 0.5629880, 0.1542950, 0.6970960, 0.3636720, 0.8959430, 0.9580330, 0.1638830, 0.9638650, 0.0403664, 0.4740620, 0.6345540, 0.2606130, 0.8029370, 0.9051410, 0.3828440, 0.2208010, 0.5651010, 0.6397810, 0.1436260, 0.4426360, 0.2803950, 0.2998880, 0.0791335, 0.2059480, 0.6069810, 0.5667200, 0.4700820, 0.3595450, 0.2252730, 0.8470000, 0.6382970, 0.4591530, 0.9537550, 0.2336280, 0.3840740, 0.7791530, 0.1905040, 0.0379216, 0.0795039, 0.6224730, 0.2131420, 0.7705720, 0.7632950, 0.1969430, 0.9052830, 0.5194640, 0.9537460, 0.9094010, 0.1706940, 0.0162099, 0.3670480, 0.6247680, 0.7822800, 0.6563370, 0.8297280, 0.0365994, 0.1534690, 0.1695770, 0.8372420, 0.5863690, 0.4421480, 0.9581610, 0.2074660, 0.9404130, 0.5156770, 0.1751960, 0.8746480, 0.8116410, 0.6343980, 0.5525990, 0.6126000, 0.9128680, 0.9037180, 0.1081180, 0.2430410, 0.2621660, 0.0548171, 0.2393530, 0.9490780, 0.2504170, 0.0771853, 0.2508970, 0.6902880, 0.6040980, 0.3622870, 0.0535081, 0.0686587, 0.2101600, 0.0907458, 0.2109090, 0.6404060, 0.3476860, 0.6944910, 0.0614566, 0.0508914, 0.6219590, 0.0488251, 0.7301400, 0.7823590, 0.1846250, 0.9812910, 0.5652960, 0.3983750, 0.1956970, 0.6458630, 0.8840490, 0.5769660, 0.1283370, 0.2979040, 0.7862870, 0.3184020, 0.8284230, 0.9035590, 0.1387210, 0.7427180, 0.1012920, 0.6461890, 0.6374320, 0.8309130, 0.2094780, 0.5971390, 0.2762440, 0.3904880, 0.1913530, 0.1954260, 0.1136790, 0.8275850, 0.6065680, 0.9592890, 0.2093050, 0.7565840, 0.5886220, 0.0783072, 0.5186390, 0.6247440, 0.7084760, 0.5537470, 0.6867080, 0.7320310, 0.9742790, 0.1631280, 0.3074160, 0.3978790, 0.2441060, 0.9211560, 0.9427770, 0.1557330, 0.0939716, 0.6561770, 0.8017070, 0.6074040, 0.7286530, 0.8264550, 0.6716160, 0.7528690, 0.6526280, 0.3964640, 0.1489860, 0.2308810, 0.3463510, 0.1519640, 0.8833840, 0.0911013, 0.9127660, 0.0389184, 0.6478400, 0.9476410, 0.6696680, 0.4743090, 0.3377090, 0.8883880, 0.9831240, 0.4802090, 0.2226000, 0.8435670, 0.6143130, 0.2817880, 0.1987060, 0.2756800, 0.6718370, 0.2704100, 0.7912680, 0.0221030, 0.5096260, 0.1372450, 0.9430530, 0.9772590, 0.8562300, 0.9656660, 0.1214440, 0.7900540, 0.9448010, 0.6546670, 0.0802318, 0.8411850, 0.8038360, 0.7777670, 0.5959040, 0.0936029, 0.9227380, 0.1135310, 0.9516650, 0.2254730, 0.4265170, 0.0696742, 0.6619350, 0.2703240, 0.1646940, 0.4126910, 0.6162690, 0.1587070, 0.3520620, 0.0298689, 0.1641180, 0.8869670, 0.5133290, 0.5606760, 0.6495700, 0.8499110, 0.2489560, 0.0272232, 0.0658381, 0.8177920, 0.3111810, 0.1596590, 0.7275860, 0.5664260, 0.3487670, 0.5039090, 0.5749390, 0.3608460, 0.3921370, 0.1024180, 0.5346650, 0.7273790, 0.9548820, 0.8175060, 0.8815920, 0.7927300, 0.6396790, 0.9801550, 0.0039532, 0.1092690, 0.9278640, 0.5746140, 0.4604150, 0.6435760, 0.7050270, 0.9683830, 0.0393886, 0.1857360, 0.6608870, 0.4605380, 0.9894990, 0.8834680, 0.6240120, 0.8934090, 0.7029980, 0.8359460, 0.3809430, 0.2062450, 0.9354910, 0.3905090, 0.2415100, 0.1506150, 0.8793510, 0.6014540, 0.7273380, 0.3160260, 0.9050160, 0.8643800, 0.2187550, 0.1895550, 0.3408190, 0.2138430, 0.9554440, 0.7446450, 0.8057730, 0.0007480, 0.5884090, 0.9320450, 0.9788700, 0.7651770, 0.4800880, 0.4909470, 0.2952700, 0.3218100, 0.7579970, 0.5694070, 0.8112590, 0.7876230, 0.8345740, 0.6259230, 0.7930130, 0.7643430, 0.1826500, 0.6887810, 0.3934710, 0.9224670, 0.3350110, 0.7139600, 0.8245460, 0.0626045, 0.6179420, 0.3326470, 0.8213810, 0.7862520, 0.3132390, 0.8836740, 0.4040760, 0.6952120, 0.2019920, 0.5085220, 0.6432880, 0.3217630, 0.0308972, 0.7565570, 0.4211240, 0.0131949, 0.3624330, 0.2708860, 0.0707916, 0.3997690, 0.7490850, 0.2423490, 0.7423600, 0.3110500, 0.7874400, 0.6439920, 0.8216780, 0.9197490, 0.8084260, 0.8770630, 0.8374480, 0.4928090, 0.6812780, 0.4958270, 0.6048640, 0.9405300, 0.5209420, 0.9461410, 0.7567610, 0.7679060, 0.3510630, 0.3719420, 0.2602230, 0.4851010, 0.3574090, 0.9240840, 0.2397680, 0.3298580, 0.4465260, 0.7666970, 0.8031800, 0.4806210, 0.8401600, 0.4932150, 0.9566480, 0.9235720, 0.2663930, 0.7974970, 0.1999000, 0.1758790, 0.9321940, 0.3201670, 0.5680990, 0.5586450, 0.7846910, 0.2438620, 0.4884790, 0.1273190, 0.2268940, 0.9825270, 0.6471090, 0.9317380, 0.7770530, 0.1431020, 0.2879080, 0.4410940, 0.3629390, 0.5319860, 0.5746750, 0.4780390, 0.2875500, 0.5514210, 0.6336410, 0.8757520, 0.0566193, 0.6524400, 0.8015120, 0.3319970, 0.0875375, 0.9028770, 0.2569820, 0.6602440, 0.6846360, 0.1931570, 0.6601510, 0.5339920, 0.9502640, 0.1829560, 0.3889620, 0.9971170, 0.4904460, 0.7848520, 0.5374680, 0.1200820, 0.7892350, 0.3970620, 0.4105070, 0.6771450, 0.5875720, 0.7336880, 0.0574303, 0.5303240, 0.2445590, 0.9443490, 0.8904020, 0.6390250, 0.3619560, 0.8266500, 0.0674818, 0.3571580, 0.7636370, 0.7685470, 0.5139750, 0.8354260, 0.1669520, 0.9379460, 0.7153450, 0.5212920, 0.9179660, 0.2712450, 0.7964090, 0.3452930, 0.4070340, 0.7370710, 0.5793780, 0.9995340, 0.7446760, 0.2363040, 0.0561258, 0.1880760, 0.8681960, 0.9400790, 0.3716920, 0.3887590, 0.8214270, 0.6420110, 0.4760180, 0.7875780, 0.7024290, 0.7755740, 0.9840510, 0.1603240, 0.7016030, 0.9026740, 0.8163780, 0.2291300, 0.4573230, 0.6498620, 0.8890870, 0.3945890, 0.7159140, 0.7975940, 0.4209690, 0.1948190, 0.7003340, 0.3677480, 0.9230850, 0.1717690, 0.4488600, 0.4043810, 0.9952960, 0.8496350, 0.4606770, 0.1002120, 0.7165120, 0.6708700, 0.2851850, 0.7324310, 0.2068220, 0.1767720, 0.7891610, 0.7320210, 0.4606250, 0.6794960, 0.1466770, 0.7657460, 0.2221640, 0.0178033, 0.6109490, 0.4956960, 0.7587780, 0.9942500, 0.9105670, 0.2693280, 0.7057770, 0.6026390, 0.3643530, 0.4193120, 0.4448910, 0.4177640, 0.8950320, 0.6667370, 0.2169620, 0.4441530, 0.2289370, 0.5174220, 0.0357793, 0.3906260, 0.3419230, 0.9172170, 0.3616600, 0.6422970, 0.9185450, 0.5705750, 0.3447180, 0.0088229, 0.5684610, 0.0100397, 0.5729230, 0.3318520, 0.8674990, 0.9931050, 0.2024440, 0.3410200, 0.5999840, 0.8546760, 0.7378130, 0.6395390, 0.7974410, 0.0319022, 0.7257180, 0.2874060, 0.6047000, 0.8955910, 0.2768590, 0.1471240, 0.2768850, 0.0622604, 0.5840070, 0.0561934, 0.2529030, 0.4694260, 0.4812150, 0.8479970, 0.3290990, 0.4851870, 0.8243810, 0.2776060, 0.3581150, 0.4834690, 0.4930710, 0.0917412, 0.0845144, 0.2188840, 0.2136950, 0.7318320, 0.5751890, 0.3305610, 0.5673700, 0.3466350, 0.3081220, 0.1295800, 0.3336710, 0.2896680, 0.1258770, 0.6128230, 0.4673290, 0.5420330, 0.2777600, 0.2004720, 0.4007360, 0.9061960, 0.2367780, 0.0635779, 0.1744970, 0.1668280, 0.0207054, 0.1895550, 0.4739310, 0.2811160, 0.2870790, 0.9346070, 0.2051150, 0.0349663, 0.6358760, 0.5394670, 0.7203070, 0.2952550, 0.2654630, 0.9802030, 0.6000470, 0.6222820, 0.3932450, 0.1008950, 0.2018130, 0.8025190, 0.6942880, 0.6448740, 0.6309640, 0.4293630, 0.9242380, 0.2566920, 0.7208310, 0.7055140, 0.6346100, 0.9811470, 0.2992960, 0.9985590, 0.9960810, 0.0087002, 0.6654140, 0.0963863, 0.1917060, 0.6426700, 0.1025770, 0.4215890, 0.2808810, 0.0167665, 0.3908970, 0.5053870, 0.3261210, 0.1995350, 0.9791030, 0.9354930, 0.4889110, 0.2520670, 0.5791210, 0.1998740, 0.5346720, 0.2728780, 0.2374600, 0.7587430, 0.4748830, 0.0052523, 0.9941600, 0.7064580, 0.9822530, 0.7476780, 0.4103290, 0.5778920, 0.4340100, 0.0440194, 0.6032060, 0.5637070, 0.1105720, 0.1515170, 0.8335130, 0.5701900, 0.4345250, 0.0657179, 0.5060150, 0.2973670, 0.4018860, 0.1950820, 0.8165790, 0.8700140, 0.7425550, 0.5313820, 0.5261480, 0.7106650, 0.5902050, 0.9514570, 0.6531750, 0.4436010, 0.8501960, 0.7745300, 0.7136690, 0.5192740, 0.1056420, 0.9074410, 0.1214610, 0.6324500, 0.4051580, 0.9777230, 0.5074190, 0.8007910, 0.1730870, 0.7570390, 0.7369090, 0.1438690, 0.1905500, 0.4660520, 0.9484070, 0.4488180, 0.6292740, 0.3441000, 0.7657860, 0.3941330, 0.8863430, 0.7340290, 0.0493191, 0.6259250, 0.5315000, 0.4721680, 0.2644180, 0.9149140, 0.6238340, 0.9919960, 0.3612810, 0.8815700, 0.8668770, 0.2125820, 0.1670860, 0.3368520, 0.5948730, 0.7963890, 0.1482670, 0.8873710, 0.5036960, 0.0313617, 0.0658449, 0.8495830, 0.8511190, 0.6914480, 0.9232690, 0.2087660, 0.1283130, 0.0910550, 0.3657740, 0.9889910, 0.3500040, 0.4745320, 0.7687570, 0.4291030, 0.1870430, 0.3664060, 0.5215910, 0.6113800, 0.4378540, 0.2493290, 0.8962560, 0.9610800, 0.2750510, 0.3055250, 0.2887760, 0.9533340, 0.3074340, 0.5237370, 0.5694600, 0.4415970, 0.1942730, 0.1059130, 0.4408260, 0.7727600, 0.0651168, 0.5501230, 0.0911351, 0.1141330, 0.5292510, 0.5326990, 0.0630471, 0.9129740, 0.0066872, 0.1326640, 0.8407100, 0.7230720, 0.2649980, 0.1925590, 0.5194330, 0.9668590, 0.2311120, 0.7283650, 0.3482210, 0.3889630, 0.2833100, 0.8447800, 0.2401950, 0.4218880, 0.9387150, 0.0025263, 0.6480120, 0.6834780, 0.1839070, 0.8378620, 0.9200110, 0.7942620, 0.1708400, 0.5348020, 0.4090720, 0.3330680, 0.3602580, 0.7075360, 0.1005620, 0.3195760, 0.4912660, 0.5946390, 0.2626710, 0.7981100, 0.6272940, 0.3476090, 0.8346990, 0.4827580, 0.3282310, 0.0987056, 0.3860400, 0.7132420, 0.4228550, 0.1204980, 0.0745314, 0.3338790, 0.4699790, 0.5063100, 0.0884488, 0.1581430, 0.4026900, 0.8763140, 0.8862410, 0.9076170, 0.6581660, 0.9217070, 0.0752826, 0.5366720, 0.0601108, 0.3512140, 0.2445370, 0.9712720, 0.5863210, 0.6800990, 0.0416432, 0.8682560, 0.9435910, 0.8797700, 0.6996800, 0.8825220, 0.4259660, 0.5834920, 0.6970860, 0.9927150, 0.1919060, 0.1573270, 0.3544910, 0.0842331, 0.1512280, 0.6375530, 0.5288450, 0.4716290, 0.7772750, 0.6119770, 0.2728070, 0.9823210, 0.5995340, 0.1109320, 0.9544510, 0.3799930, 0.4938070, 0.4469910, 0.3593660, 0.4491400, 0.5164730, 0.5553610, 0.8751630, 0.5059840, 0.9484300, 0.9729110, 0.3143850, 0.6781020, 0.7776020, 0.8965090, 0.2291660, 0.8256450, 0.6814280, 0.2404050, 0.6902070, 0.3692700, 0.6851190, 0.0350788, 0.3185510, 0.3648830, 0.4334940, 0.6320970, 0.4355490, 0.0191081, 0.6847580, 0.7946160, 0.7860570, 0.3720360, 0.8627480, 0.4283790, 0.0832822, 0.2941540, 0.8150520, 0.9061870, 0.7756530, 0.6545660, 0.8794370, 0.4802560, 0.4596130, 0.8941020, 0.4883160, 0.8479060, 0.5374710, 0.9719620, 0.2561120, 0.4904100, 0.8619420, 0.7367310, 0.6701930, 0.0655039, 0.4144210, 0.0659039, 0.5244620, 0.5794410, 0.2513870, 0.9415480, 0.3294540, 0.8732670, 0.9302620, 0.3635740, 0.7783660, 0.5531730, 0.7952030, 0.2828690, 0.4433060, 0.1653840, 0.6146930, 0.0297614, 0.8927450, 0.7269480, 0.4547570, 0.0965830, 0.4592100, 0.1617840, 0.0729463, 0.0502157, 0.8518920, 0.8084450, 0.5771590, 0.3435940, 0.9214080, 0.0448326, 0.5212360, 0.4611200, 0.0561864, 0.6028330, 0.8618160, 0.1525980, 0.1532170, 0.3198590, 0.9551610, 0.4539760, 0.5176480, 0.0825359, 0.6349380, 0.3494150, 0.4514320, 0.5748300, 0.4032290, 0.8533680, 0.0046974, 0.0998581, 0.8289600, 0.7843870, 0.0163287, 0.3615860, 0.0039164, 0.3414110, 0.9752580, 0.4431780, 0.9814760, 0.9319510, 0.4670430, 0.1941480, 0.7544260, 0.4769630, 0.0605473, 0.1495700, 0.1351880, 0.2389690, 0.7767920, 0.4620700, 0.0839400, 0.7791500, 0.9013870, 0.4346180, 0.0194434, 0.1108420, 0.2433440, 0.2236820, 0.2814690, 0.5872330, 0.9138110, 0.0588877, 0.7518610, 0.3118460, 0.0626417, 0.7941540, 0.8278480, 0.5524520, 0.7176670, 0.6756500, 0.8050770, 0.9052880, 0.0302903, 0.3153700, 0.5394880, 0.4674020, 0.9505300, 0.1398640, 0.8063700, 0.1271010, 0.6325780, 0.0804024, 0.8462380, 0.4896780, 0.7189560, 0.3634970, 0.9884420, 0.3695290, 0.3271360, 0.8505420, 0.6352760, 0.2610650, 0.7561170, 0.1735160, 0.8133560, 0.3108930, 0.2419100, 0.5314590, 0.1909310, 0.5459960, 0.5894850, 0.8460650, 0.8136500, 0.4256290, 0.5384500, 0.7218600, 0.5115490, 0.3795100, 0.5703850, 0.8168150, 0.4792140, 0.6115120, 0.8238100, 0.1250150, 0.9944810, 0.2605130, 0.2772430, 0.1680330, 0.6830380, 0.9240380, 0.9712460, 0.2255810, 0.2121740, 0.1603070, 0.4178910, 0.2600720, 0.6710360, 0.7117600, 0.3075860, 0.3039980, 0.9560810, 0.2004160, 0.7370170, 0.1207890, 0.0553623, 0.2329920, 0.3399640, 0.0433382, 0.0162401, 0.0589458, 0.0231145, 0.4469360, 0.7397640, 0.7408910, 0.4416140, 0.0964111, 0.7014520, 0.0925169, 0.7352000, 0.4348590, 0.4394570, 0.8883580, 0.6960280, 0.6612080, 0.3694020, 0.1086570, 0.2864540, 0.0385367, 0.1676570, 0.3426510, 0.5392900, 0.4753730, 0.9427260, 0.0666164, 0.0060144, 0.2943750, 0.0733364, 0.6951760, 0.3501700, 0.4683150, 0.0259394, 0.7216030, 0.2277790, 0.7162830, 0.8442900, 0.8654280, 0.9499720, 0.0423316, 0.0717323, 0.8904640, 0.9684530, 0.9136820, 0.9698760, 0.7841690, 0.9841490, 0.5646770, 0.4478400, 0.0981987, 0.1966330, 0.7967610, 0.0071249, 0.9885710, 0.0024369, 0.7790160, 0.5188000, 0.1136310, 0.1756170, 0.0430181, 0.1328680, 0.4137150, 0.8751130, 0.0689622, 0.6862480, 0.7868110, 0.9013580, 0.6115040, 0.5822240, 0.2009900, 0.5872860, 0.1089340, 0.3855130, 0.3625430, 0.2997770, 0.1837570, 0.1409040, 0.2231560, 0.2191020, 0.2520120, 0.1454860, 0.1735300, 0.8400810, 0.9507130, 0.0539245, 0.3751640, 0.2744020, 0.3096190, 0.4343820, 0.5698470, 0.7054990, 0.2045640, 0.1768770, 0.1828840, 0.3547910, 0.0662873, 0.6594180, 0.6941040, 0.9594500, 0.9123850, 0.1035170, 0.3758250, 0.7977830, 0.5142650, 0.0024239, 0.2020720, 0.0735932, 0.9041270, 0.3662850, 0.2963760, 0.1325770, 0.9444680, 0.7904760, 0.8382900, 0.9921950, 0.3833490, 0.3159580, 0.5282360, 0.3876680, 0.6392590, 0.7430920, 0.1039730, 0.9673910, 0.2554960, 0.6481680, 0.1049840, 0.3674880, 0.1139570, 0.4768500, 0.4355060, 0.0592776, 0.1887360, 0.8100500, 0.4528890, 0.1597240, 0.5918600, 0.6393070, 0.6097040, 0.4035540, 0.0851091, 0.6914690, 0.2095460, 0.1260500, 0.3405380, 0.8710980, 0.3940060, 0.7720870, 0.1727030, 0.5582670, 0.3483940, 0.1145390, 0.3456310, 0.1570970, 0.0928358, 0.3278720, 0.2632950, 0.7620350, 0.6706560, 0.5709520, 0.3561110, 0.9300780, 0.4151060, 0.5250000, 0.3279380, 0.5897250, 0.7323890, 0.7401830, 0.9169780, 0.5351890, 0.3366010, 0.5802670, 0.8904040, 0.7862170, 0.3118910, 0.3270140, 0.9201680, 0.2429740, 0.2890520, 0.0771307, 0.6645350, 0.8208590, 0.8633320, 0.8162160, 0.7815550, 0.1771610, 0.5533450, 0.0787490, 0.0204303, 0.0768594, 0.7665890, 0.4871160, 0.3050870, 0.8787000, 0.1290380, 0.1602660, 0.7638680, 0.8317800, 0.6762830, 0.9443300, 0.6466050, 0.8423210, 0.7777100, 0.3792210, 0.2463250, 0.5809390, 0.1663090, 0.4397100, 0.4683730, 0.5911540, 0.4770800, 0.7290410, 0.1099830, 0.3974400, 0.5282260, 0.3629260, 0.9026290, 0.2892660, 0.8472230, 0.2000270, 0.5265300, 0.0564947, 0.0574168, 0.2360760, 0.5302580, 0.1591540, 0.3618050, 0.4050650, 0.6995990, 0.6508000, 0.9989620, 0.3410080, 0.3195430, 0.1158160, 0.5904700, 0.9270210, 0.2231930, 0.9210870, 0.9496840, 0.4003810, 0.7588190, 0.1155920, 0.3354380, 0.8575360, 0.6882830, 0.0681853, 0.6331940, 0.0750319, 0.6614400, 0.5083260, 0.2754800, 0.5477760, 0.5508860, 0.3245280, 0.5464370, 0.6696060, 0.3952440, 0.7673130, 0.7595970, 0.6254450, 0.2789630, 0.6532600, 0.7102920, 0.3075640, 0.0513375, 0.2701740, 0.6946930, 0.2925420, 0.1629300, 0.8388410, 0.4095540, 0.1903630, 0.2685820, 0.0392356, 0.9521940, 0.6481580, 0.3684180, 0.1385390, 0.4791630, 0.5838310, 0.3144750, 0.3516660, 0.7721720, 0.7356800, 0.3754270, 0.3884370, 0.9872780, 0.4548270, 0.2850480, 0.2904990, 0.9574660, 0.6955300, 0.1848090, 0.7058440, 0.7416190, 0.1300200, 0.3817730, 0.3203860, 0.3609440, 0.8501330, 0.6907580, 0.8286910, 0.4813810, 0.0749817, 0.3077210, 0.3970540, 0.4698750, 0.1338400, 0.4730260, 0.9340890, 0.4533110, 0.3646770, 0.8830980, 0.8485740, 0.0863663, 0.4932600, 0.7954040, 0.1960600, 0.2616420, 0.3769780, 0.4313720, 0.3028150, 0.8882370, 0.5822670, 0.3571430, 0.2004270, 0.1451980, 0.5170870, 0.7258000, 0.8528810, 0.1383860, 0.4410170, 0.1844290, 0.9891350, 0.6078740, 0.2462780, 0.1269620, 0.5358040, 0.4410170, 0.0428544, 0.9427390, 0.7339070, 0.9725020, 0.1708040, 0.1366130, 0.9074580, 0.2776990, 0.6366700, 0.4384880, 0.0068678, 0.4195770, 0.3159400, 0.1386780, 0.1044970, 0.2296250, 0.3393130, 0.2735060, 0.3183510, 0.4017860, 0.7151800, 0.0296360, 0.7332910, 0.3450080, 0.7444050, 0.4561240, 0.9601760, 0.0707048, 0.2308440, 0.0492430, 0.1405300, 0.3172180, 0.3149380, 0.8271580, 0.6126690, 0.1618240, 0.8052220, 0.3264740, 0.4473340, 0.3951830, 0.3940910, 0.9492130, 0.8348680, 0.6984040, 0.3107890, 0.0126802, 0.0088530, 0.7083510, 0.4807190, 0.1134100, 0.3268790, 0.1269500, 0.2964410, 0.5201670, 0.2734200, 0.3217140, 0.7010220, 0.3769510, 0.9139570, 0.0843911, 0.9644940, 0.7926710, 0.6230750, 0.0102056, 0.3375270, 0.0654856, 0.0542729, 0.0302635, 0.3626260, 0.7222170, 0.4384830, 0.6726310, 0.5214250, 0.9435120, 0.0304840, 0.1230060, 0.6207940, 0.0102451, 0.1802880, 0.8633710, 0.8161870, 0.5643690, 0.4846060, 0.7639460, 0.0828837, 0.3162840, 0.2504220, 0.3950340, 0.7656090, 0.9662330, 0.2994610, 0.0526907, 0.3513080, 0.3683570, 0.8223170, 0.7196030, 0.1753020, 0.8198890, 0.2320590, 0.2307440, 0.0009750, 0.0666662, 0.5239170, 0.4040550, 0.4325950, 0.2882900, 0.6646980, 0.3885980, 0.3715890, 0.5437530, 0.8599410, 0.3173910, 0.5540770, 0.3875790, 0.4346350, 0.2289280, 0.8087830, 0.0207723, 0.8852230, 0.0684584, 0.6903380, 0.9554720, 0.0848232, 0.2542280, 0.3555830, 0.2909900, 0.6144600, 0.6168310, 0.0737309, 0.0619436, 0.0506739, 0.2477320, 0.4722440, 0.1299770, 0.1487830, 0.6236970, 0.0579531, 0.1445550, 0.4488910, 0.4514590, 0.4091420, 0.6326580, 0.3707500, 0.7387270, 0.2192830, 0.4790330, 0.0911552, 0.8694200, 0.1550700, 0.3067940, 0.0322670, 0.4857370, 0.8598650, 0.4245730, 0.7693190, 0.6234420, 0.5625180, 0.8584470, 0.4573250, 0.6211330, 0.3247190, 0.8264670, 0.3885440, 0.4098780, 0.1073970, 0.8469500, 0.5078570, 0.6592330, 0.9518900, 0.2845090, 0.5965510, 0.9433370, 0.6272170, 0.6839970, 0.1935130, 0.4654030, 0.2086220, 0.9374500, 0.5165380, 0.9964920, 0.0998501, 0.1474570, 0.3833380, 0.8860190, 0.5060720, 0.8003350, 0.4281920, 0.2639110, 0.5684220, 0.5599450, 0.4608390, 0.2999280, 0.2511000, 0.1952740, 0.5767900, 0.4197040, 0.7319830, 0.7969620, 0.8268370, 0.7538950, 0.6176600, 0.9906700, 0.6158360, 0.4198110, 0.1851820, 0.1478700, 0.0347870, 0.6212160, 0.3240200, 0.0648480, 0.8489010, 0.0270243, 0.6690370, 0.5566390, 0.8729700, 0.0015362, 0.0216633, 0.3433100, 0.9006970, 0.2731130, 0.3572780, 0.7268220, 0.6089010, 0.6865130, 0.7404200, 0.3319570, 0.0779955, 0.3676940, 0.7150960, 0.1862250, 0.3673610, 0.6986840, 0.6336200, 0.0593625, 0.5916590, 0.5576550, 0.9654090, 0.5903040, 0.6512010, 0.5733590, 0.1999740, 0.6341510, 0.5038560, 0.4794600, 0.7479880, 0.4040200, 0.0337409, 0.0931086, 0.7824130, 0.2229310, 0.8594180, 0.1160440, 0.6677170, 0.5452230, 0.9600140, 0.0570182, 0.3857730, 0.8902140, 0.2911260, 0.0232105, 0.1410780, 0.5273030, 0.7108280, 0.8352910, 0.8026120, 0.6001630, 0.4121860, 0.6045540, 0.1988380, 0.5826900, 0.9250200, 0.3355500, 0.3904160, 0.5858300, 0.0714631, 0.9590400, 0.9450710, 0.4868570, 0.6252130, 0.4813510, 0.2741180, 0.5537640, 0.3400170, 0.6423660, 0.4796390, 0.2755010, 0.7665570, 0.7529830, 0.1329100, 0.9959910, 0.5350300, 0.2843520, 0.2784080, 0.6284320, 0.3236140, 0.8120230, 0.1806490, 0.1025950, 0.8866330, 0.0394051, 0.9077550, 0.3016320, 0.9860890, 0.7222920, 0.4564790, 0.6819880, 0.2364200, 0.8525970, 0.3955510, 0.7125130, 0.7747120, 0.4665530, 0.7272320, 0.9748170, 0.2443110, 0.8988360, 0.0490816, 0.9441900, 0.4422270, 0.0684266, 0.2119730, 0.4139380, 0.2333700, 0.2860880, 0.5255900, 0.7635780, 0.4088560, 0.8064340, 0.1876680, 0.6323830, 0.0672180, 0.0814072, 0.3392150, 0.8681310, 0.8343420, 0.5182250, 0.8419780, 0.9534060, 0.4751980, 0.9377420, 0.7694170, 0.2021090, 0.8249290, 0.3481410, 0.9389250, 0.9445160, 0.7694980, 0.1353250, 0.3237050, 0.7531350, 0.3009690, 0.9710990, 0.0341473, 0.9982290, 0.7851200, 0.6639170, 0.2608920, 0.6232060, 0.9628880, 0.5096470, 0.6487000, 0.3266630, 0.6648820, 0.9563700, 0.4206770, 0.2175470, 0.4218540, 0.7942700, 0.4070510, 0.8778300, 0.9146820, 0.6724740, 0.9332790, 0.4009190, 0.8208290, 0.4960760, 0.1140190, 0.7695680, 0.8265730, 0.3757980, 0.7662280, 0.8981470, 0.8008770, 0.8702440, 0.9228170, 0.4418140, 0.6161940, 0.6373120, 0.4259030, 0.8820910, 0.4498130, 0.3928210, 0.7477430, 0.2613450, 0.0942952, 0.0976953, 0.3769440, 0.3474160, 0.7813960, 0.4034120, 0.5897320, 0.9223230, 0.8051450, 0.3585150, 0.1913430, 0.9935880, 0.7230370, 0.7126210, 0.9206480, 0.5129450, 0.4394070, 0.5797020, 0.7060260, 0.3540790, 0.3598930, 0.9039160, 0.9607940, 0.6882930, 0.1673420, 0.2877110, 0.3095770, 0.3439260, 0.0875487, 0.1333950, 0.9379430, 0.4687460, 0.2216650, 0.7747970, 0.7067680, 0.5523990, 0.7048900, 0.4637820, 0.0001386, 0.6055620, 0.3206280, 0.7280750, 0.1837640, 0.9218940, 0.0965211, 0.6701450, 0.4794090, 0.8093920, 0.8619310, 0.2963690, 0.2637170, 0.8975740, 0.6621640, 0.3307770, 0.7026500, 0.7212560, 0.6681050, 0.3785880, 0.6151790, 0.4889010, 0.8948480, 0.6733950, 0.4556570, 0.4428000, 0.6941410, 0.6428600, 0.3467390, 0.9828380, 0.2674400, 0.8175840, 0.5636450, 0.2238630, 0.3636550, 0.1108930, 0.6650930, 0.7789150, 0.1745810, 0.6629230, 0.1413410, 0.3767320, 0.4487020, 0.0200910, 0.6615400, 0.6407690, 0.3443290, 0.6969680, 0.0999750, 0.1398460, 0.2296490, 0.0278118, 0.1612550, 0.2166160, 0.5188670, 0.5524930, 0.2788270, 0.4958190, 0.7062660, 0.3488530, 0.7972640, 0.7939650, 0.0636304, 0.4670420, 0.9674380, 0.8073900, 0.8539100, 0.1079130, 0.4827580, 0.5161260, 0.9320800, 0.3942780, 0.7538780, 0.9546090, 0.3119540, 0.5008830, 0.0735425, 0.7881350, 0.1691890, 0.3123000, 0.8595270, 0.9789450, 0.6705450, 0.2845310, 0.3433620, 0.2682540, 0.2409520, 0.4825400, 0.3806880, 0.5894350, 0.0915371, 0.5332460, 0.8774250, 0.5256980, 0.7879000, 0.3066830, 0.1772740, 0.4367750, 0.3010750, 0.8643750, 0.7113360, 0.2442030, 0.6562480, 0.1644080, 0.9489210, 0.6994980, 0.5921770, 0.0604606, 0.0131991, 0.8832000, 0.8163590, 0.4971010, 0.8590040, 0.8066100, 0.3491790, 0.3040990, 0.2183840, 0.8971270, 0.8918740, 0.5885550, 0.9401470, 0.0033195, 0.9060990, 0.6317710, 0.5955040, 0.6108410, 0.5339710, 0.9674360, 0.7455060, 0.6176140, 0.2036100, 0.2381850, 0.3112120, 0.6144070, 0.6281520, 0.3981860, 0.6260780, 0.4136490, 0.1227850, 0.4034710, 0.3630750, 0.6833200, 0.5693070, 0.3359460, 0.9633190, 0.4639970, 0.9402680, 0.2069180, 0.6116540, 0.7619620, 0.7646540, 0.5254700, 0.0404121, 0.3353330, 0.8312750, 0.2487040, 0.5429460, 0.9061120, 0.4696000, 0.4443040, 0.1058940, 0.2542650, 0.9738240, 0.1915140, 0.0492553, 0.5023770, 0.3008560, 0.6554960, 0.4814340, 0.3137970, 0.5373700, 0.0328781, 0.1932270, 0.6258780, 0.9916570, 0.2327890, 0.8760970, 0.4994190, 0.9349470, 0.5467850, 0.2101650, 0.4217340, 0.9147500, 0.3175440, 0.5781340, 0.3133670, 0.2820600, 0.9631280, 0.3449490, 0.8392260, 0.3194900, 0.3595670, 0.5612670, 0.5762080, 0.4846160, 0.8079530, 0.9011240, 0.1061410, 0.1134750, 0.6868120, 0.1837650, 0.7002940, 0.4321850, 0.6428730, 0.4252050, 0.0664025, 0.0174651, 0.3855020, 0.3762960, 0.8977370, 0.7679690, 0.7124530, 0.8600600, 0.2524310, 0.9166990, 0.0221280, 0.3680150, 0.8943120, 0.7778890, 0.8316680, 0.8329700, 0.2935290, 0.5068260, 0.7280200, 0.8658080, 0.8197720, 0.8795710, 0.6509920, 0.5598090, 0.2159320, 0.8500670, 0.3613170, 0.2927360, 0.4817610, 0.0630102, 0.1925050, 0.8770410, 0.9520730, 0.1187570, 0.9962350, 0.1876010, 0.1774890, 0.2742410, 0.3051670, 0.8830760, 0.4622380, 0.1200800, 0.5333700, 0.9001160, 0.8985870, 0.6005960, 0.1788550, 0.5882080, 0.2858760, 0.9919180, 0.1729120, 0.9775310, 0.5499110, 0.7912770, 0.5005610, 0.9262410, 0.3138320, 0.4270020, 0.1918440, 0.5562320, 0.4610820, 0.5797890, 0.2745240, 0.8522120, 0.1974100, 0.8523930, 0.0024974, 0.0006961, 0.2027320, 0.9025600, 0.9325750, 0.9610840, 0.8261050, 0.3119160, 0.8163000, 0.9900800, 0.9083130, 0.7046770, 0.2874830, 0.9041310, 0.1425820, 0.9059440, 0.4467050, 0.1764980, 0.8633980, 0.0375420, 0.7692250, 0.4633820, 0.9768730, 0.8282710, 0.5012960, 0.7764970, 0.7019540, 0.2580910, 0.9728840, 0.3709770, 0.0589938, 0.9215440, 0.8718060, 0.2874240, 0.8728610, 0.9723370, 0.0907140, 0.3218360, 0.1701850, 0.0589483, 0.1306280, 0.6259550, 0.1164550, 0.8546460, 0.2065380, 0.7420150, 0.1659220, 0.2006350, 0.4742780, 0.5107250, 0.3346220, 0.3400860, 0.8766490, 0.5493340, 0.0682539, 0.2763480, 0.3269260, 0.1349170, 0.6181080, 0.8953400, 0.4118610, 0.0335518, 0.3520980, 0.8091160, 0.9352540, 0.7027610, 0.9181150, 0.5972430, 0.3985020, 0.2200400, 0.4603600, 0.6227340, 0.4260680, 0.9008130, 0.5815010, 0.8956670, 0.1757580, 0.2773330, 0.0374825, 0.2892200, 0.0516494, 0.2079110, 0.5028910, 0.7497240, 0.9124400, 0.2215000, 0.5866900, 0.7813060, 0.6117080, 0.9450980, 0.5259350, 0.3590160, 0.9361330, 0.0787932, 0.9212970, 0.9889590, 0.3362330, 0.4232230, 0.4976790, 0.9250090, 0.6537010, 0.5638170, 0.4241980, 0.3882220, 0.2293450, 0.2657450, 0.6322070, 0.3710700, 0.5050260, 0.9332500, 0.9681630, 0.2674990, 0.4730080, 0.9193210, 0.7715980, 0.7341790, 0.2236620, 0.6468210, 0.4894000, 0.9020330, 0.3361520, 0.4754650, 0.5042510, 0.7142850, 0.0938567, 0.7007110, 0.2662740, 0.3929630, 0.9382840, 0.0504546, 0.1255380, 0.8863360, 0.1013010, 0.3671150, 0.7426240, 0.1475920, 0.2551200, 0.9735000, 0.6462370, 0.1756350, 0.0370002, 0.1338590, 0.6362810, 0.3633870, 0.4430670, 0.8717280, 0.6242760, 0.2015920, 0.7253660, 0.7926460, 0.1498460, 0.4172290, 0.5359100, 0.7188330, 0.4042640, 0.7323010, 0.2844980, 0.8809850, 0.8935600, 0.6661480, 0.0828788, 0.8445560, 0.9821710, 0.7662310, 0.7553750, 0.6834470, 0.9234290, 0.4605180, 0.5916770, 0.5015180, 0.0528082, 0.8809030, 0.9568320, 0.2108070, 0.2659540, 0.1347990, 0.6480910, 0.7385520, 0.1532470, 0.0212134, 0.0680201, 0.6134310, 0.8163480, 0.1501310, 0.4200550, 0.3483940, 0.7181380, 0.3124760, 0.9460500, 0.0097909, 0.2213540, 0.9934480, 0.1957270, 0.8727360, 0.5290780, 0.8529550, 0.9592700, 0.5187290, 0.7889360, 0.3343410, 0.8668540, 0.9658020, 0.9958750, 0.3264090, 0.7296440, 0.3942870, 0.7271610, 0.0543889, 0.3825630, 0.5108650, 0.8206090, 0.2571590, 0.5861630, 0.5138340, 0.6992930, 0.5720210, 0.4346030, 0.6622970, 0.0877279, 0.2301620, 0.2333550, 0.1619080, 0.5818180, 0.3852310, 0.2514820, 0.4733210, 0.8610510, 0.5895720, 0.0548549, 0.9732100, 0.2725510, 0.3677380, 0.9294190, 0.0036511, 0.3771990, 0.7026410, 0.0718129, 0.5127010, 0.7418490, 0.7180140, 0.6279430, 0.4486320, 0.8492420, 0.8314120, 0.5963990, 0.2906780, 0.8033110, 0.6324880, 0.0077729, 0.2257170, 0.4314710, 0.5963080, 0.9803380, 0.2432500, 0.0864019, 0.3561750, 0.7368110, 0.3657440, 0.8471070, 0.2972330, 0.8720180, 0.7512410, 0.4001670, 0.2422590, 0.2819230, 0.7059180, 0.5723560, 0.2421110, 0.8662340, 0.7741940, 0.5154000, 0.0346658, 0.1155590, 0.8172400, 0.1662520, 0.0593847, 0.5228370, 0.1481520, 0.9849670, 0.5010640, 0.8607690, 0.3634500, 0.6171530, 0.3734360, 0.0022691, 0.5939120, 0.9071030, 0.9612430, 0.1748730, 0.2469880, 0.1362940, 0.8733300, 0.1104200, 0.4960530, 0.0417473, 0.6525950, 0.0923936, 0.6169090, 0.1406250, 0.3860670, 0.6272510, 0.5786950, 0.0473607, 0.5650900, 0.7110260, 0.5071060, 0.5286910, 0.1306270, 0.6224750, 0.4934870, 0.7303940, 0.8899770, 0.8891110, 0.7703980, 0.2790870, 0.2604850, 0.7789410, 0.8598370, 0.9067990, 0.6750910, 0.4551580, 0.9160570, 0.6037520, 0.0111074, 0.3477360, 0.5254250, 0.8757220, 0.5419490, 0.0530215, 0.1058750, 0.5032910, 0.5874140, 0.3879720, 0.0663841, 0.9420470, 0.3554800, 0.8843090, 0.0453011, 0.3301000, 0.3833590, 0.0669687, 0.1549260, 0.9783380, 0.5359390, 0.9257200, 0.9949090, 0.7538790, 0.0093842, 0.9357840, 0.1784190, 0.8268900, 0.9596760, 0.9585460, 0.0516299, 0.2063460, 0.4183420, 0.7159140, 0.2374010, 0.7278990, 0.4339140, 0.4617030, 0.4940750, 0.9779170, 0.2130810, 0.5447380, 0.3152310, 0.5479190, 0.3601150, 0.1493320, 0.6749930, 0.1713640, 0.9682380, 0.3473420, 0.1523220, 0.8713770, 0.4229210, 0.2460770, 0.5205790, 0.0914422, 0.0578432, 0.8235290, 0.6495690, 0.7865480, 0.3213320, 0.7431450, 0.5296800, 0.7829140, 0.7619780, 0.1877800, 0.8663120, 0.0667691, 0.2050110, 0.4549960, 0.1880180, 0.1047300, 0.6187870, 0.7394030, 0.7489810, 0.0511937, 0.7199790, 0.5387970, 0.9591980, 0.6547020, 0.8140170, 0.1957450, 0.4846330, 0.0078575, 0.4523440, 0.8081720, 0.8136840, 0.1827970, 0.4834200, 0.7307250, 0.3900280, 0.6609710, 0.4059410, 0.1636720, 0.9367010, 0.0955379, 0.0717113, 0.1629700, 0.3270330, 0.1532440, 0.3080230, 0.1166930, 0.7817760, 0.4756170, 0.0533785, 0.4412740, 0.8305770, 0.1611590, 0.2136480, 0.6920160, 0.2686980, 0.6790690, 0.9774880, 0.0089960, 0.6550350, 0.0708997, 0.1464170, 0.7315860, 0.7485200, 0.0304747, 0.1124730, 0.2657890, 0.3746260, 0.5361730, 0.4615750, 0.5047510, 0.4420640, 0.3603920, 0.9634750, 0.8789890, 0.8423020, 0.7547960, 0.9565690, 0.9324280, 0.2414240, 0.6253170, 0.2635360, 0.6270470, 0.4143270, 0.6082950, 0.8778260, 0.9548300, 0.5080980, 0.1003660, 0.1155040, 0.7313500, 0.6814420, 0.1451900, 0.8142300, 0.9184420, 0.8447860, 0.6725680, 0.3297630, 0.3308630, 0.3465490, 0.8720970, 0.5967160, 0.8960170, 0.6734850, 0.1127590, 0.5568260, 0.4371690, 0.2918950, 0.4056250, 0.7461460, 0.7697250, 0.5139090, 0.3129460, 0.7003900, 0.4558270, 0.8319770, 0.8393560, 0.9011830, 0.7996600, 0.4344270, 0.3249680, 0.2207150, 0.1631060, 0.9712280, 0.0990465, 0.5285840, 0.2583210, 0.2897410, 0.4745330, 0.5440050, 0.4719180, 0.4622720, 0.6253370, 0.5325510, 0.3923890, 0.5985840, 0.2110950, 0.3718380, 0.0856160, 0.7085480, 0.1829720, 0.7844340, 0.0290660, 0.9417690, 0.9160300, 0.4391930, 0.8095320, 0.1416440, 0.9856590, 0.4285560, 0.4011480, 0.2069700, 0.3037520, 0.5826960, 0.0024956, 0.3966000, 0.3897520, 0.4705290, 0.2559700, 0.9359660, 0.5962500, 0.1693930, 0.0402567, 0.3393180, 0.2856010, 0.2676420, 0.1093300, 0.0838898, 0.2218030, 0.2109480, 0.3898130, 0.7658890, 0.2306220, 0.5664320, 0.2596390, 0.9569150, 0.3707750, 0.8027720, 0.6694960, 0.7457370, 0.1732590, 0.3440540, 0.7715840, 0.2548460, 0.3067980, 0.0003238, 0.4731130, 0.9983230, 0.7680440, 0.1849260, 0.6324050, 0.3472910, 0.1697510, 0.0546478, 0.4085470, 0.1774010, 0.1924250, 0.5909490, 0.6641900, 0.2927680, 0.8992840, 0.7646230, 0.8283350, 0.5249060, 0.4315810, 0.7720560, 0.3747050, 0.9559240, 0.6682550, 0.8484990, 0.6187120, 0.4186620, 0.9363960, 0.5633350, 0.7185060, 0.2553740, 0.0329907, 0.5456020, 0.5492600, 0.4623610, 0.8619250, 0.9961200, 0.3005570, 0.7132860, 0.3647770, 0.2906470, 0.1039760, 0.6250440, 0.4369140, 0.2526440, 0.0992564, 0.1899470, 0.5417550, 0.5830800, 0.8533680, 0.9418040, 0.4217160, 0.8744250, 0.0607349, 0.6978790, 0.3764140, 0.9413990, 0.7734640, 0.2643890, 0.9583290, 0.6611440, 0.6403120, 0.0353324, 0.5371780, 0.3652280, 0.1902520, 0.8807930, 0.1766420, 0.4007250, 0.1177600, 0.4407840, 0.0901711, 0.1578890, 0.6433300, 0.1838700, 0.0758178, 0.3192560, 0.5646950, 0.0502260, 0.4522310, 0.5532320, 0.2244600, 0.1710650, 0.0495389, 0.3593680, 0.2518970, 0.4188800, 0.6062270, 0.6240550, 0.4676180, 0.2518580, 0.0012189, 0.5617040, 0.2027020, 0.9864150, 0.5674150, 0.4449820, 0.6539280, 0.4378980, 0.9183270, 0.5938680, 0.9430030, 0.4058160, 0.5353540, 0.4560570, 0.3793890, 0.8373440, 0.4444310, 0.4505100, 0.8610350, 0.7897230, 0.2233990, 0.0424224, 0.8020500, 0.8777670, 0.9401130, 0.7924670, 0.8498040, 0.1051550, 0.6400970, 0.0307505, 0.0601553, 0.9647230, 0.3393400, 0.6537830, 0.8697460, 0.9631810, 0.2592620, 0.2553710, 0.8942490, 0.2812120, 0.5190500, 0.1817390, 0.6607980, 0.8108570, 0.6408110, 0.0444925, 0.8241110, 0.9938310, 0.9236590, 0.5857450, 0.3986910, 0.7670430, 0.8376140, 0.7271520, 0.0501445, 0.9464650, 0.0199312, 0.3620340, 0.6133800, 0.9662530, 0.7142280, 0.1006200, 0.9124210, 0.8843340, 0.1045480, 0.6174070, 0.7200030, 0.9500720, 0.2830860, 0.3333780, 0.5336130, 0.1815110, 0.4644800, 0.2328810, 0.7253280, 0.9062500, 0.8289350, 0.7726700, 0.3750340, 0.5742110, 0.2171940, 0.7721860, 0.2454010, 0.6764960, 0.7237040, 0.0413954, 0.8737190, 0.0090614, 0.4008110, 0.9691330, 0.6768640, 0.2977790, 0.0071465, 0.9155320, 0.5946420, 0.3580620, 0.5178350, 0.8899650, 0.0815958, 0.7236850, 0.2612000, 0.2397920, 0.6129340, 0.2056470, 0.5981810, 0.7347470, 0.2485940, 0.4356840, 0.5572200, 0.9706010, 0.5484210, 0.2096100, 0.6707270, 0.0109817, 0.0818821, 0.3301210, 0.2843140, 0.2433160, 0.6264200, 0.8244470, 0.2645130, 0.4895610, 0.7259680, 0.8268620, 0.4423220, 0.7106960, 0.1565580, 0.5959930, 0.1538350, 0.5242770, 0.0047548, 0.3541530, 0.3395620, 0.5375730, 0.0974282, 0.3263080, 0.9925460, 0.2579380, 0.1131200, 0.8244700, 0.9155700, 0.4597220, 0.0821045, 0.7342580, 0.8647960, 0.0160573, 0.3583770, 0.2581610, 0.2991910, 0.5266640, 0.8059820, 0.0803884, 0.6776490, 0.0938045, 0.3680130, 0.5077910, 0.9212480, 0.6176690, 0.2040430, 0.3260280, 0.9278270, 0.1868950, 0.1965720, 0.4419170, 0.0847753, 0.3402740, 0.6757100, 0.1455500, 0.1749830, 0.1673350, 0.8361290, 0.4691830, 0.3914590, 0.6123430, 0.3510230, 0.2774110, 0.8653970, 0.8511180, 0.4182600, 0.7105210, 0.2445470, 0.4384060, 0.5230470, 0.9942290, 0.8995440, 0.0228073, 0.6343740, 0.6742740, 0.0907487, 0.6998580, 0.0218377, 0.1981120, 0.4202180, 0.5980260, 0.4977360, 0.1433570, 0.5351630, 0.7158880, 0.5156800, 0.0523013, 0.5321800, 0.5802370, 0.6793780, 0.7157290, 0.5951100, 0.1582540, 0.2689960, 0.8534340, 0.5980600, 0.0908210, 0.5305670, 0.6101610, 0.3550180, 0.7293340, 0.1673120, 0.2909590, 0.3549100, 0.8523150, 0.5739280, 0.2163990, 0.0127750, 0.7206290, 0.0053457, 0.0724694, 0.7324950, 0.5894530, 0.7467340, 0.3641990, 0.7851690, 0.8282770, 0.1173800, 0.2985040, 0.3806570, 0.1791530, 0.4900070, 0.2829660, 0.5055070, 0.0202066, 0.4320820, 0.5706960, 0.0035709, 0.3769520, 0.6725210, 0.1282760, 0.0760981, 0.8019060, 0.4100780, 0.6105030, 0.1005100, 0.4823550, 0.0161053, 0.3974840, 0.2736390, 0.0253331, 0.0072673, 0.0637050, 0.1368880, 0.4252520, 0.2302370, 0.4925650, 0.9160790, 0.9618720, 0.1379090, 0.0425270, 0.5389340, 0.2687710, 0.9132700, 0.7723480, 0.2597950, 0.4343910, 0.4502980, 0.5182510, 0.4943750, 0.6457220, 0.8571750, 0.4311110, 0.4396000, 0.2301780, 0.1029060, 0.0256695, 0.4841630, 0.8929220, 0.7436050, 0.9953460, 0.9289490, 0.6164260, 0.3546360, 0.3108620, 0.5398870, 0.3120590, 0.6017240, 0.6361570, 0.1443940, 0.0584834, 0.7399090, 0.5282060, 0.5513710, 0.5756990, 0.0259969, 0.0443242, 0.7764370, 0.3380990, 0.6706520, 0.0356107, 0.6151100, 0.4849920, 0.0706852, 0.2098120, 0.4902490, 0.0855852, 0.3332330, 0.5975590, 0.2977430, 0.0200496, 0.2028170, 0.2127770, 0.4581560, 0.7184450, 0.7984770, 0.3259280, 0.4691010, 0.7522880, 0.8885330, 0.3365730, 0.3902780, 0.9908910, 0.1703780, 0.8384890, 0.4614580, 0.1500000, 0.2709910, 0.9029520, 0.6592840, 0.3327940, 0.3289450, 0.6114300, 0.7594430, 0.5841100, 0.4412080, 0.8116720, 0.8758330, 0.6188660, 0.4027660, 0.3192280, 0.2439730, 0.1567360, 0.2889310, 0.7280740, 0.1786450, 0.8893870, 0.1783890, 0.0838219, 0.5656790, 0.5489680, 0.3070030, 0.8751690, 0.5730230, 0.6742930, 0.4106970, 0.2341910, 0.4046830, 0.2670590, 0.0324075, 0.1161570, 0.9678710, 0.2582750, 0.8645460, 0.5587290, 0.4950660, 0.9339760, 0.5479900, 0.1925870, 0.5930200, 0.4897500, 0.5390550, 0.4434050, 0.7356910, 0.4745130, 0.1050480, 0.6729250, 0.5660740, 0.8772940, 0.9048160, 0.2968760, 0.0643319, 0.8936430, 0.4555810, 0.6225750, 0.2594860, 0.4995000, 0.1003750, 0.4690550, 0.4820370, 0.9226450, 0.2516970, 0.6565590, 0.5254910, 0.0926267, 0.9886030, 0.6590720, 0.7085290, 0.7147330, 0.3360470, 0.3332140, 0.9601870, 0.0069907, 0.0348025, 0.1579980, 0.3252610, 0.3309120, 0.3237850, 0.9881770, 0.7097750, 0.6949760, 0.7337540, 0.8968930, 0.5261660, 0.5701380, 0.0250271, 0.4184500, 0.0214821, 0.7216230, 0.4594510, 0.2044610, 0.7075100, 0.3111800, 0.7304590, 0.9543730, 0.7195960, 0.7313480, 0.8796320, 0.3790800, 0.1565950, 0.6091980, 0.9096660, 0.7455540, 0.3317170, 0.6039200, 0.7733980, 0.8635640, 0.3375020, 0.1361310, 0.1781290, 0.4426440, 0.4984650, 0.3445600, 0.3301680, 0.8557720, 0.0880057, 0.0403901, 0.1922000, 0.4553240, 0.2761110, 0.6244410, 0.0114162, 0.4635500, 0.2591640, 0.9963120, 0.7624700, 0.2709880, 0.0276698, 0.8620020, 0.1092410, 0.6638910, 0.5755700, 0.8146280, 0.2559840, 0.8204990, 0.4207000, 0.0580771, 0.3114700, 0.8554740, 0.8772000, 0.9930380, 0.4643220, 0.3333920, 0.0976139, 0.9823300, 0.8630300, 0.1547530, 0.5247820, 0.2075420, 0.5207120, 0.9728030, 0.9029940, 0.8913280, 0.1812880, 0.1337980, 0.7492310, 0.6058830, 0.5119300, 0.4333000, 0.9689010, 0.7329540, 0.8573860, 0.7231940, 0.0154615, 0.8827040, 0.0848824, 0.7659870, 0.5181200, 0.8653550, 0.3904370, 0.9982260, 0.9134130, 0.4848260, 0.7119200, 0.8970430, 0.8749700, 0.6848810, 0.0314156, 0.6322670, 0.8870390, 0.6811750, 0.9930570, 0.8962530, 0.9084940, 0.9606850, 0.9426750, 0.1024160, 0.6078760, 0.8874980, 0.2336900, 0.5789410, 0.8469470, 0.5382620, 0.3076860, 0.1622740, 0.7908390, 0.5478850, 0.0074982, 0.1393000, 0.1967000, 0.9414250, 0.1554360, 0.3249590, 0.0681518, 0.4186290, 0.2798510, 0.9088190, 0.6176240, 0.3745830, 0.7498310, 0.2727400, 0.5689210, 0.8883190, 0.1982250, 0.5256770, 0.7688970, 0.1355970, 0.8553930, 0.5692950, 0.9917050, 0.5181890, 0.6113460, 0.9986970, 0.1131820, 0.3589420, 0.7572760, 0.2902920, 0.4995920, 0.1810820, 0.2428710, 0.4049250, 0.5442410, 0.5644210, 0.6810680, 0.3664090, 0.5961210, 0.7776620, 0.4050110, 0.5217140, 0.0340909, 0.9247400, 0.2637600, 0.7616900, 0.0551694, 0.7747900, 0.3113600, 0.7369170, 0.8736280, 0.1625280, 0.5357520, 0.9271730, 0.6349980, 0.1812960, 0.7310380, 0.2540920, 0.5254400, 0.2891800, 0.3141040, 0.5248890, 0.4100550, 0.6928150, 0.4045800, 0.5631480, 0.7292900, 0.6141060, 0.6060650, 0.9242190, 0.1037890, 0.6590520, 0.2338940, 0.8145120, 0.5136650, 0.1684450, 0.2007090, 0.7484220, 0.0305673, 0.5167320, 0.8717620, 0.5690800, 0.6185680, 0.3372100, 0.6494520, 0.7515400, 0.7174890, 0.0249133, 0.3186230, 0.2162050, 0.0409259, 0.0601466, 0.6771410, 0.4885290, 0.2729080, 0.5661630, 0.3831620, 0.5738140, 0.8095240, 0.3658450, 0.4530570, 0.5977460, 0.8041630, 0.1974830, 0.9427680, 0.3770020, 0.9222360, 0.1685510, 0.3863980, 0.1230200, 0.0183627, 0.6510800, 0.9088140, 0.9822220, 0.9027950, 0.9600390, 0.8009030, 0.4659010, 0.1663310, 0.8600090, 0.7572800, 0.9764800, 0.8871200, 0.5434080, 0.4994160, 0.2219280, 0.2940720, 0.9719490, 0.0165047, 0.7264370, 0.1281530, 0.5368300, 0.3691380, 0.1864550, 0.1725320, 0.3480760, 0.0914221, 0.0776030, 0.0023043, 0.3344920, 0.9664520, 0.3841780, 0.7056600, 0.3974460, 0.3370360, 0.1294580, 0.7394910, 0.5357270, 0.5666060, 0.1500650, 0.2588630, 0.5364610, 0.6235360, 0.8374790, 0.0958546, 0.3801050, 0.4183080, 0.9161340, 0.0136536, 0.4302320, 0.1527350, 0.7171980, 0.8582410, 0.4376430, 0.7668950, 0.4621670, 0.7355360, 0.2258220, 0.8476170, 0.4971430, 0.9881620, 0.4503270, 0.4465670, 0.9050660, 0.1445830, 0.6000090, 0.9902140, 0.1707710, 0.5320190, 0.7520090, 0.8771970, 0.9884290, 0.7141420, 0.6179510, 0.4405730, 0.4932660, 0.4422960, 0.4547730, 0.7252740, 0.7664500, 0.5309030, 0.9488010, 0.0869481, 0.5622070, 0.0195833, 0.2675420, 0.2745610, 0.1383210, 0.4846280, 0.8927100, 0.8176050, 0.2144190, 0.6828000, 0.2540670, 0.5224060, 0.0135314, 0.4735180, 0.3808070, 0.4526040, 0.3482530, 0.4635750, 0.6193150, 0.9482300, 0.5527020, 0.6345270, 0.0216383, 0.4935260, 0.8633430, 0.6118090, 0.6941700, 0.4628460, 0.6642820, 0.4643370, 0.1036510, 0.0242418, 0.8645300, 0.1312120, 0.5102550, 0.9548340, 0.2499810, 0.6043190, 0.1609000, 0.7258140, 0.4226090, 0.1377820, 0.9265960, 0.8423330, 0.1310310, 0.7547910, 0.3573180, 0.2222850, 0.7929040, 0.8325540, 0.4367260, 0.2045350, 0.6457520, 0.8444090, 0.2895320, 0.2699780, 0.2761050, 0.0660376, 0.1721480, 0.3142790, 0.5002560, 0.7821120, 0.0700579, 0.7714690, 0.9481140, 0.5594110, 0.1978680, 0.5371920, 0.3928500, 0.4615130, 0.9445430, 0.1663770, 0.8057640, 0.5897780, 0.3080400, 0.7770960, 0.4871410, 0.7652240, 0.9775540, 0.4133820, 0.2742410, 0.7410340, 0.2130860, 0.7988240, 0.1737100, 0.7436430, 0.2783580, 0.3076870, 0.4745790, 0.0722817, 0.9263740, 0.4892950, 0.7581780, 0.2112770, 0.3835910, 0.8030800, 0.8297430, 0.0463752, 0.2127000, 0.6711740, 0.8283130, 0.9823200, 0.1450920, 0.4061250, 0.9345060, 0.5248640, 0.7989460, 0.9174790, 0.5440380, 0.1940340, 0.5840390, 0.3918120, 0.8600260, 0.0587082, 0.9149280, 0.3049890, 0.5375710, 0.6322110, 0.6863370, 0.7344020, 0.0989952, 0.7733210, 0.5287400, 0.9102210, 0.7433950, 0.8308370, 0.1903530, 0.8950350, 0.3920020, 0.6627800, 0.3013540, 0.2825490, 0.2272900, 0.7356000, 0.3094150, 0.9101850, 0.9463290, 0.3562720, 0.4934630, 0.0005187, 0.5335230, 0.6432830, 0.6094800, 0.3149030, 0.6312720, 0.0940048, 0.4526870, 0.5219890, 0.7572680, 0.5362680, 0.5149900, 0.9475470, 0.3243510, 0.7910730, 0.6991110, 0.0360273, 0.6289980, 0.2311060, 0.3788960, 0.0062391, 0.7125650, 0.8747400, 0.7982170, 0.0094399, 0.6301180, 0.8987230, 0.2833800, 0.5034670, 0.7703450, 0.9643320, 0.7936620, 0.7531800, 0.4140370, 0.5858380, 0.3897460, 0.4266630, 0.8352940, 0.9043590, 0.6668250, 0.4301370, 0.4773520, 0.8021280, 0.1783620, 0.9816450, 0.0730970, 0.4630230, 0.3629130, 0.0786986, 0.6409540, 0.3771250, 0.3578130, 0.4065660, 0.0185690, 0.4150400, 0.8956890, 0.4676550, 0.4594950, 0.9577480, 0.9981870, 0.5126880, 0.4123320, 0.1823470, 0.7432640, 0.7331480, 0.8901730, 0.2665720, 0.7866210, 0.9414620, 0.3072330, 0.3026490, 0.4843740, 0.6102030, 0.2469010, 0.3244000, 0.5693430, 0.3480600, 0.8188900, 0.6980710, 0.0481705, 0.9102870, 0.0695032, 0.1155790, 0.5442800, 0.7861920, 0.2989000, 0.7819170, 0.7747330, 0.8502620, 0.9800000, 0.1166620, 0.3208180, 0.5116350, 0.7910540, 0.6718070, 0.5068380, 0.1193890, 0.0736078, 0.8646390, 0.9183870, 0.6149600, 0.5557840, 0.4239430, 0.9193810, 0.1735640, 0.5348810, 0.8228160, 0.2316740, 0.5126240, 0.5905510, 0.0853193, 0.5783950, 0.9491470, 0.9998980, 0.7194660, 0.2451690, 0.3105400, 0.3357960, 0.8017460, 0.8127340, 0.4966750, 0.8626540, 0.7094790, 0.4148590, 0.1654690, 0.4073200, 0.8951010, 0.5906870, 0.9212200, 0.1512040, 0.7597590, 0.2744650, 0.4755930, 0.7955140, 0.2122870, 0.9040790, 0.7670230, 0.6787680, 0.5908490, 0.8472270, 0.5567180, 0.0873732, 0.1769740, 0.3691200, 0.5354710, 0.3878140, 0.2945970, 0.4365070, 0.3925090, 0.0078837, 0.9021630, 0.8284600, 0.0151838, 0.2811740, 0.3280840, 0.7527680, 0.7168800, 0.6982450, 0.5900050, 0.4938300, 0.6805900, 0.2356230, 0.5285860, 0.1181550, 0.2773630, 0.2388330, 0.7684550, 0.3799860, 0.9340350, 0.5054200, 0.0540806, 0.2294260, 0.4397380, 0.8134060, 0.9521210, 0.5940880, 0.6645860, 0.4690770, 0.1409730, 0.9357190, 0.5624810, 0.8260940, 0.8375040, 0.8363240, 0.7512800, 0.9490100, 0.5833220, 0.1486950, 0.4907950, 0.2277100, 0.4499650, 0.4562630, 0.4960970, 0.9260570, 0.2659150, 0.3642800, 0.5012000, 0.3160210, 0.2535010, 0.9906480, 0.8231630, 0.5106300, 0.3910180, 0.5319040, 0.7282450, 0.5413670, 0.4343370, 0.8778990, 0.0975537, 0.7412890, 0.9671770, 0.1491490, 0.7007880, 0.4442230, 0.3066960, 0.0718324, 0.8100520, 0.4136610, 0.0030411, 0.3370360, 0.0397904, 0.5254270, 0.8828770, 0.7068000, 0.8501920, 0.5079440, 0.3621770, 0.7479760, 0.4684880, 0.0043925, 0.7286860, 0.9165170, 0.1840930, 0.4618780, 0.4011380, 0.9638560, 0.8745200, 0.0051356, 0.3045260, 0.7877700, 0.3461920, 0.0174010, 0.7779840, 0.0016535, 0.9922780, 0.9744140, 0.1800580, 0.9245780, 0.8403070, 0.5984160, 0.1174480, 0.5240780, 0.4061810, 0.2763930, 0.2672750, 0.7638970, 0.8751270, 0.4298790, 0.9409380, 0.7270830, 0.0211485, 0.5503260, 0.3136720, 0.6808910, 0.8119840, 0.1177510, 0.5076830, 0.7131660, 0.6556200, 0.2661770, 0.6880450, 0.5621630, 0.9822020, 0.4524760, 0.1895070, 0.0667989, 0.5449060, 0.8987100, 0.2486450, 0.5361830, 0.9286720, 0.5823800, 0.5329270, 0.2416630, 0.3337280, 0.8804640, 0.2920970, 0.2221870, 0.1269980, 0.4326750, 0.9839490, 0.7000790, 0.8569930, 0.9822500, 0.2741500, 0.3667860, 0.2142810, 0.2825040, 0.4558520, 0.5359620, 0.2508530, 0.0787864, 0.1308850, 0.1714450, 0.9158270, 0.6301900, 0.8561430, 0.6159730, 0.9949980, 0.4695180, 0.2664800, 0.7043870, 0.3264800, 0.2312520, 0.0632448, 0.3033320, 0.8415130, 0.5875460, 0.5734360, 0.6381020, 0.4771240, 0.1085200, 0.1458640, 0.0377676, 0.9750260, 0.2055950, 0.9921700, 0.2910150, 0.6428800, 0.2709700, 0.0598429, 0.9604680, 0.9350690, 0.5355650, 0.1003950, 0.9497030, 0.2540900, 0.6603800, 0.6506630, 0.4520170, 0.6966040, 0.0638942, 0.4140540, 0.5133920, 0.9531330, 0.7537070, 0.6831440, 0.9992970, 0.4494180, 0.3006380, 0.3213390, 0.8170490, 0.8068840, 0.6173210, 0.0417506, 0.6987030, 0.3715980, 0.9367940, 0.9649680, 0.8811170, 0.1653460, 0.1167730, 0.2898480, 0.1112970, 0.9923190, 0.3739940, 0.8491110, 0.2870310, 0.1175710, 0.7639780, 0.6604900, 0.3224550, 0.8858520, 0.1113700, 0.9634260, 0.4587320, 0.1999030, 0.3015260, 0.1947090, 0.0462241, 0.1127090, 0.5378300, 0.2994570, 0.5500020, 0.2442480, 0.3989670, 0.8836610, 0.7286360, 0.2075520, 0.9628240, 0.6678590, 0.3159080, 0.0411929, 0.2818580, 0.3176670, 0.6449800, 0.7959400, 0.9225710, 0.3618700, 0.8995950, 0.0417054, 0.7882670, 0.0004433, 0.5383730, 0.7936580, 0.5275780, 0.6911100, 0.9644300, 0.8114310, 0.8594630, 0.0617257, 0.5788910, 0.1122410, 0.2681800, 0.0592394, 0.5408230, 0.6751380, 0.7267580, 0.1242070, 0.4932910, 0.1196910, 0.4380720, 0.9342230, 0.9139790, 0.4980680, 0.0615753, 0.5486800, 0.2285380, 0.3806550, 0.3614360, 0.0429798, 0.5719130, 0.2552300, 0.3377100, 0.9463610, 0.7317140, 0.9222130, 0.5536420, 0.6077390, 0.5599410, 0.2961530, 0.7512360, 0.3961330, 0.1668130, 0.0730276, 0.0700529, 0.7419080, 0.1117550, 0.5357420, 0.7695900, 0.4314500, 0.1614220, 0.3938980, 0.2287700, 0.8416040, 0.7516130, 0.0899907, 0.1854410, 0.5999180, 0.4215310, 0.9725610, 0.2604660, 0.0998870, 0.3631430, 0.9784870, 0.9366010, 0.5276840, 0.0364264, 0.3183800, 0.5618170, 0.0467328, 0.4978460, 0.9486470, 0.7625830, 0.9343970, 0.9876870, 0.5028560, 0.5077880, 0.4970880, 0.7196690, 0.1896270, 0.5949990, 0.4888960, 0.6280760, 0.1540590, 0.5703400, 0.7596190, 0.0225962, 0.5157950, 0.5056380, 0.1348590, 0.6997570, 0.3025660, 0.6949890, 0.1962220, 0.3782960, 0.8100160, 0.4308820, 0.1235110, 0.3473370, 0.3142550, 0.7156110, 0.3919070, 0.8803100, 0.9317070, 0.2612940, 0.4131270, 0.4782280, 0.3421240, 0.7158140, 0.3904900, 0.1608350, 0.8673980, 0.8828840, 0.2231460, 0.0641421, 0.3735490, 0.1359440, 0.5514800, 0.7710900, 0.9350650, 0.6544490, 0.9566230, 0.3897140, 0.2533640, 0.3637430, 0.4210230, 0.4035720, 0.2349210, 0.3681060, 0.0305224, 0.5857020, 0.6365590, 0.8856950, 0.0337834, 0.2227210, 0.5543520, 0.0077415, 0.6267630, 0.0170009, 0.8288250, 0.3295770, 0.8455910, 0.9095340, 0.4085840, 0.8262230, 0.1449170, 0.8033000, 0.9716560, 0.7324500, 0.7342300, 0.8379450, 0.2176470, 0.4662490, 0.3624990, 0.0419045, 0.2291830, 0.1741820, 0.1664470, 0.0838837, 0.2727260, 0.8151690, 0.3714170, 0.4401950, 0.8741000, 0.6742780, 0.1078350, 0.3924890, 0.2479830, 0.4786750, 0.9188080, 0.9596940, 0.5793330, 0.9912720, 0.4733070, 0.3599020, 0.4678490, 0.7272820, 0.8889630, 0.4785690, 0.1177970, 0.8760770, 0.4033940, 0.2720690, 0.4581960, 0.6006420, 0.3882640, 0.7433050, 0.6997690, 0.1923960, 0.9984310, 0.4339680, 0.7593220, 0.4646780, 0.6086660, 0.2171980, 0.2971050, 0.6154880, 0.7708660, 0.1566680, 0.2944820, 0.1941930, 0.7956380, 0.9027760, 0.8563050, 0.4063570, 0.9464450, 0.8324810, 0.7013420, 0.7177190, 0.3199220, 0.9950850, 0.5761380, 0.4630820, 0.1894050, 0.4911810, 0.2169740, 0.1430340, 0.0402711, 0.7434120, 0.5974760, 0.3122370, 0.1978560, 0.8798000, 0.7556350, 0.4281340, 0.1648690, 0.6696080, 0.7420140, 0.8328450, 0.2912480, 0.9545550, 0.8690450, 0.0452972, 0.1436010, 0.8134570, 0.7349720, 0.2077930, 0.7234740, 0.4910440, 0.3767420, 0.0544776, 0.1218140, 0.0599685, 0.3440290, 0.6186680, 0.0663865, 0.4225870, 0.7456330, 0.1247630, 0.3399370, 0.8859980, 0.7412500, 0.8580130, 0.1308200, 0.6074740, 0.3059820, 0.5814630, 0.2059170, 0.2526660, 0.8143560, 0.4909230, 0.3027940, 0.3668490, 0.1025600, 0.7459650, 0.5507830, 0.5591130, 0.2375190, 0.3581320, 0.3695950, 0.2344820, 0.0912443, 0.3592580, 0.0187052, 0.9294860, 0.4014110, 0.3817770, 0.9889830, 0.6249610, 0.8856510, 0.5221700, 0.9189630, 0.1218850, 0.4382350, 0.8691780, 0.0064826, 0.5198100, 0.2675690, 0.9653360, 0.2263600, 0.1040520, 0.8339600, 0.3852230, 0.6773180, 0.3730370, 0.3647490, 0.2570730, 0.1053370, 0.3207380, 0.2641030, 0.3367080, 0.8877830, 0.6023830, 0.9677250, 0.3623060, 0.9376910, 0.2638820, 0.1514710, 0.2945850, 0.3922430, 0.5301470, 0.6060070, 0.4341610, 0.8805340, 0.1854540, 0.7414420, 0.7659610, 0.9420370, 0.6829690, 0.3188870, 0.4849390, 0.8749420, 0.6501340, 0.7202770, 0.6090110, 0.6242730, 0.4979820, 0.5642550, 0.3740310, 0.6973250, 0.9539430, 0.1555020, 0.5973890, 0.6545630, 0.2553850, 0.6170700, 0.4601030, 0.0335217, 0.3415600, 0.9890800, 0.7403400, 0.3247960, 0.8030100, 0.2966310, 0.7444400, 0.5311720, 0.5708600, 0.2728320, 0.4384620, 0.4015550, 0.0024445, 0.0392649, 0.3229990, 0.3625140, 0.6019470, 0.4596190, 0.2420390, 0.4812400, 0.3053410, 0.4507060, 0.3871950, 0.7685030, 0.6306700, 0.0168539, 0.8671040, 0.7492640, 0.9877620, 0.5749190, 0.3674620, 0.8406670, 0.5376940, 0.5064210, 0.1889820, 0.7727690, 0.4596230, 0.8957800, 0.4695030, 0.8989310, 0.8974950, 0.6895470, 0.0519178, 0.1982410, 0.0626402, 0.9297640, 0.6101510, 0.6423960, 0.0032043, 0.7472680, 0.4242730, 0.9048560, 0.8844720, 0.0604422, 0.9778630, 0.4684240, 0.2946340, 0.3682620, 0.4402670, 0.9750390, 0.8337670, 0.1486090, 0.4379930, 0.3592010, 0.6964630, 0.2186540, 0.5628930, 0.0037381, 0.7257110, 0.1976960, 0.8385980, 0.3708300, 0.6197680, 0.6343490, 0.9308630, 0.8824760, 0.6047040, 0.2237730, 0.0793241, 0.4677930, 0.8675740, 0.1409660, 0.5727580, 0.4314280, 0.0543695, 0.7333830, 0.1904710, 0.9475010, 0.0989259, 0.0988213, 0.7939320, 0.1475610, 0.5290390, 0.0201558, 0.1956900, 0.4543100, 0.2053280, 0.3956490, 0.6509090, 0.7880770, 0.8117550, 0.1516190, 0.6345580, 0.0487502, 0.6644640, 0.3865620, 0.4620270, 0.6169000, 0.0384687, 0.1473360, 0.0826269, 0.6994410, 0.2210550, 0.3441640, 0.1724820, 0.8689200, 0.7556590, 0.0412911, 0.0651409, 0.7376130, 0.5646610, 0.5609210, 0.9101370, 0.4666680, 0.2941060, 0.1440080, 0.4440620, 0.1269690, 0.8351840, 0.3068690, 0.7240800, 0.5504600, 0.9044340, 0.6738580, 0.8881400, 0.9132600, 0.7159500, 0.5408510, 0.0369161, 0.9450790, 0.5424510, 0.4897320, 0.2983280, 0.2908340, 0.8027280, 0.6376650, 0.0712580, 0.8803090, 0.9991860, 0.5175180, 0.8503080, 0.8649970, 0.6570920, 0.6484870, 0.7903660, 0.0397087, 0.9664510, 0.0870565, 0.3020020, 0.1871240, 0.1176910, 0.5105040, 0.0676704, 0.9401090, 0.8865230, 0.7741790, 0.9909560, 0.9061850, 0.5173470, 0.8430390, 0.7428790, 0.5844070, 0.5961480, 0.7588540, 0.3358040, 0.1775800, 0.6391320, 0.3264280, 0.4242720, 0.3062870, 0.8316000, 0.9007990, 0.3141810, 0.1550170, 0.3290870, 0.6620310, 0.4331500, 0.2648160, 0.2937830, 0.6596260, 0.9484250, 0.0375481, 0.6549510, 0.6210430, 0.9560830, 0.5819250, 0.4250800, 0.7143750, 0.2017800, 0.7955300, 0.9362430, 0.5071000, 0.5443270, 0.5347480, 0.6261680, 0.0972368, 0.3546320, 0.1373120, 0.5499720, 0.6402230, 0.9026530, 0.0012045, 0.1914520, 0.1227430, 0.8224560, 0.6404900, 0.5945910, 0.4064260, 0.2430280, 0.9340120, 0.3040000, 0.9139090, 0.7048310, 0.9918600, 0.4874820, 0.6993670, 0.2704350, 0.7457750, 0.4943470, 0.1966020, 0.6312080, 0.0931066, 0.4072620, 0.5752020, 0.2626390, 0.6013370, 0.3265020, 0.8081910, 0.1590620, 0.1711220, 0.2939890, 0.0316500, 0.2386310, 0.2823400, 0.1865770, 0.9178740, 0.6794850, 0.8619730, 0.5047150, 0.4990880, 0.4520530, 0.0028955, 0.0852474, 0.1909280, 0.4111060, 0.6199760, 0.8566350, 0.3495190, 0.3509750, 0.5351310, 0.7414230, 0.8141300, 0.0206768, 0.6344640, 0.4722060, 0.0984854, 0.6343700, 0.5448980, 0.9106550, 0.2764860, 0.3243000, 0.2665380, 0.0080301, 0.8373590, 0.6746320, 0.2861970, 0.0911595, 0.8335480, 0.3069380, 0.4228520, 0.3444830, 0.3545670, 0.5995330, 0.1760300, 0.5067410, 0.9453060, 0.2711960, 0.5441250, 0.5321280, 0.6601010, 0.6272220, 0.0672056, 0.8211770, 0.3290290, 0.0692197, 0.3176690, 0.7999330, 0.4604860, 0.0028980, 0.0373186, 0.3527360, 0.1988920, 0.0452814, 0.9843620, 0.3285540, 0.7438540, 0.4431400, 0.3584920, 0.5603060, 0.4905960, 0.5618620, 0.5097940, 0.9971630, 0.2997880, 0.9715230, 0.2401170, 0.4096750, 0.3268580, 0.5848430, 0.7877330, 0.0760634, 0.3742170, 0.6147080, 0.3314530, 0.4019820, 0.4435540, 0.9064760, 0.8761090, 0.5485600, 0.1870670, 0.5978760, 0.8799200, 0.6743300, 0.0427488, 0.6251640, 0.4482060, 0.0448379, 0.9733010, 0.2224720, 0.3109590, 0.6731880, 0.4299710, 0.0215786, 0.1353610, 0.6212930, 0.6692560, 0.4374750, 0.0123820, 0.1074780, 0.6542230, 0.9752190, 0.6458720, 0.0390652, 0.4134720, 0.2849790, 0.8541260, 0.3554060, 0.1770360, 0.0699990, 0.0634352, 0.1327490, 0.4402640, 0.8084060, 0.0902772, 0.8245190, 0.8577930, 0.5626560, 0.7611000, 0.1138690, 0.5134110, 0.6018090, 0.8278180, 0.4717740, 0.4303520, 0.1229760, 0.3049900, 0.5500180, 0.0669764, 0.3255830, 0.6350890, 0.5394830, 0.4737140, 0.7111920, 0.8883630, 0.5631540, 0.1353890, 0.8980930, 0.3361600, 0.7932720, 0.0337875, 0.1341460, 0.7656960, 0.3643290, 0.1466390, 0.1988820, 0.5817040, 0.6303410, 0.5732990, 0.4255370, 0.3834180, 0.9679010, 0.5244700, 0.7439480, 0.4475340, 0.0670205, 0.8435910, 0.9483030, 0.2162870, 0.5948790, 0.0039552, 0.1232780, 0.7067860, 0.7359960, 0.7363870, 0.2686590, 0.0289755, 0.3161860, 0.2867070, 0.5335890, 0.9667520, 0.1538160, 0.5456930, 0.8291870, 0.8495270, 0.3901870, 0.6166290, 0.2209090, 0.8647230, 0.1610190, 0.9125900, 0.1516040, 0.0955601, 0.0792363, 0.9020920, 0.7305350, 0.8047730, 0.5410210, 0.8966650, 0.3400780, 0.1849670, 0.3218230, 0.9303800, 0.7139450, 0.1344170, 0.8918990, 0.6152040, 0.6401580, 0.8196130, 0.9600210, 0.9728880, 0.1365200, 0.8911380, 0.7823180, 0.3862450, 0.1761860, 0.3253140, 0.0872713, 0.3834100, 0.0369643, 0.2039210, 0.8565160, 0.5791910, 0.9919040, 0.6747210, 0.0096948, 0.7276770, 0.2415890, 0.9274430, 0.9716850, 0.4994580, 0.2835880, 0.8567230, 0.8173080, 0.8515630, 0.3090280, 0.0821761, 0.6398990, 0.3408460, 0.7153100, 0.5585360, 0.8960310, 0.4551170, 0.5870590, 0.1525850, 0.9075810, 0.5291600, 0.7775180, 0.2159010, 0.5846560, 0.2689810, 0.3328290, 0.5557470, 0.4510470, 0.6715900, 0.1500360, 0.2221600, 0.5039300, 0.8110400, 0.1196280, 0.0942700, 0.9033450, 0.6898230, 0.9436510, 0.3049760, 0.1876950, 0.4100760, 0.5635850, 0.5513770, 0.7940950, 0.0136660, 0.9791380, 0.3292120, 0.5375630, 0.1308980, 0.4966890, 0.1546710, 0.4334720, 0.0160265, 0.5623520, 0.4156330, 0.7007080, 0.1097310, 0.7464650, 0.8428070, 0.0621063, 0.8183530, 0.9893080, 0.7099470, 0.7046730, 0.1391950, 0.8883360, 0.1087010, 0.6790060, 0.0823787, 0.1626870, 0.2441890, 0.0529455, 0.9314130, 0.3880940, 0.1449510, 0.3031740, 0.4311070, 0.9628660, 0.2030580, 0.2436490, 0.2155600, 0.3753810, 0.0178499, 0.1720910, 0.4844460, 0.7527240, 0.3297210, 0.5273290, 0.6991120, 0.2258710, 0.6614640, 0.0086986, 0.3899350, 0.5650440, 0.2221610, 0.9089180, 0.6026240, 0.5107920, 0.4774350, 0.9247400, 0.9468840, 0.4713010, 0.4965020, 0.8787610, 0.4669250, 0.4517880, 0.9037410, 0.0206357, 0.3953940, 0.2462590, 0.4051840, 0.2724210, 0.6063500, 0.2170090, 0.5168700, 0.1615770, 0.3170050, 0.5190330, 0.7041910, 0.8901820, 0.4692120, 0.7489060, 0.3358750, 0.2997940, 0.3036240, 0.0905017, 0.4839280, 0.6216920, 0.2420910, 0.5541790, 0.3144300, 0.8733750, 0.3091780, 0.6650900, 0.4576420, 0.1042750, 0.8936040, 0.7073040, 0.7155140, 0.3699210, 0.1683520, 0.0484401, 0.0483841, 0.8863750, 0.5324510, 0.7353110, 0.4408200, 0.0351107, 0.7962440, 0.8816530, 0.3998840, 0.8926510, 0.8437140, 0.1657220, 0.3357860, 0.9846290, 0.4991830, 0.8500860, 0.0756198, 0.7862540, 0.1231910, 0.3039750, 0.6141510, 0.3751220, 0.8915750, 0.5672660, 0.9232150, 0.7960180, 0.6100990, 0.2307640, 0.5731070, 0.6706860, 0.2127560, 0.5910310, 0.8459420, 0.9478400, 0.0908068, 0.4303520, 0.4835510, 0.1412000, 0.2882480, 0.6246290, 0.2758090, 0.3990210, 0.7825520, 0.2102950, 0.7408600, 0.5979070, 0.9505490, 0.1140640, 0.3897990, 0.3434600, 0.0592354, 0.8339900, 0.0814588, 0.6133160, 0.8669630, 0.6743060, 0.0231881, 0.0883666, 0.9532300, 0.0518525, 0.8400010, 0.2759240, 0.0934482, 0.7233820, 0.0479577, 0.7227280, 0.8111380, 0.9719970, 0.2955890, 0.4912890, 0.8238620, 0.2848500, 0.4389530, 0.5167980, 0.4013150, 0.7291720, 0.3584180, 0.3639010, 0.2246360, 0.7605350, 0.0259420, 0.9165320, 0.5800760, 0.1539810, 0.6905470, 0.7751440, 0.7179130, 0.8741430, 0.4136490, 0.7197880, 0.5878370, 0.3857030, 0.4859670, 0.5123450, 0.5608270, 0.8098110, 0.0387506, 0.8773230, 0.2074620, 0.8256110, 0.2284540, 0.9117710, 0.9470370, 0.9031020, 0.0364356, 0.1976430, 0.6688070, 0.2674890, 0.8539990, 0.2876060, 0.6649640, 0.8858640, 0.8529130, 0.7710610, 0.1337160, 0.8617310, 0.7391170, 0.0822483, 0.8497550, 0.6006740, 0.8368570, 0.9394980, 0.7488030, 0.8906760, 0.8665110, 0.6547380, 0.9053700, 0.4197350, 0.2225820, 0.3732460, 0.9144620, 0.5202180, 0.7844290, 0.5099860, 0.2350040, 0.4852920, 0.4720820, 0.1232210, 0.0833054, 0.0488025, 0.3455510, 0.9534430, 0.6433150, 0.6617240, 0.0852565, 0.5459270, 0.4885740, 0.5200150, 0.3168200, 0.8029190, 0.6962460, 0.8672860, 0.3338090, 0.7728610, 0.5038710, 0.3975260, 0.1813740, 0.0902579, 0.3874620, 0.6263970, 0.0264613, 0.2340600, 0.6264390, 0.1224770, 0.1335930, 0.5836650, 0.4052620, 0.8117560, 0.2027510, 0.2691860, 0.0295594, 0.6742860, 0.6137060, 0.2514080, 0.3794730, 0.8963420, 0.9776610, 0.3295560, 0.4095360, 0.1816500, 0.0200408, 0.4240610, 0.8988300, 0.8943810, 0.0920199, 0.7846430, 0.8666540, 0.0418388, 0.7787890, 0.6800390, 0.6086980, 0.6324600, 0.0091383, 0.1961890, 0.5570530, 0.0028572, 0.5427000, 0.6450190, 0.5846410, 0.0544814, 0.6814330, 0.5978470, 0.2933170, 0.5845300, 0.6575420, 0.4092960, 0.7001570, 0.1970640, 0.4239610, 0.9683580, 0.7807400, 0.6443410, 0.6843790, 0.8239920, 0.0034094, 0.5179130, 0.6167180, 0.8349450, 0.0262065, 0.6250130, 0.5402080, 0.7493600, 0.2912220, 0.8062860, 0.3381020, 0.7262510, 0.6295960, 0.1573000, 0.2969910, 0.9370460, 0.0766866, 0.4330000, 0.4915780, 0.0519360, 0.9134140, 0.2647260, 0.9362930, 0.3898520, 0.9979800, 0.0579981, 0.7890710, 0.0612952, 0.1398480, 0.0152750, 0.2053210, 0.8117840, 0.8082860, 0.6238910, 0.7132130, 0.5937320, 0.4643290, 0.3189960, 0.0407491, 0.4427510, 0.5214100, 0.8587440, 0.8459910, 0.2693280, 0.3352130, 0.6866950, 0.7231760, 0.7831280, 0.9439010, 0.3344300, 0.3385050, 0.9921810, 0.3704820, 0.2802240, 0.4824030, 0.9098390, 0.2612860, 0.6226420, 0.1868340, 0.7595330, 0.9439510, 0.6746930, 0.3982990, 0.8541430, 0.1658010, 0.7662290, 0.9610170, 0.9731030, 0.4671270, 0.1576410, 0.7550270, 0.3320910, 0.4889900, 0.0600297, 0.1275100, 0.1963450, 0.8529950, 0.2959630, 0.9180480, 0.3051800, 0.2269410, 0.7022040, 0.4465870, 0.4989400, 0.4554260, 0.6726690, 0.8548300, 0.2937150, 0.8293640, 0.4262880, 0.8172600, 0.7922630, 0.9866650, 0.3016760, 0.9264370, 0.3236690, 0.8124450, 0.7407120, 0.6364450, 0.0322428, 0.0813220, 0.4215590, 0.8963150, 0.4130180, 0.5504300, 0.6873990, 0.3681140, 0.0583083, 0.0424623, 0.3648620, 0.7940910, 0.8549650, 0.8319310, 0.6591180, 0.8853890, 0.0425124, 0.8090140, 0.1630900, 0.7784660, 0.2859480, 0.8052380, 0.7158860, 0.6522150, 0.1091890, 0.5486910, 0.2272950, 0.5347150, 0.4794890, 0.3925520, 0.5301890, 0.8723730, 0.5531870, 0.4002130, 0.9561430, 0.9637880, 0.5996080, 0.4254720, 0.3503220, 0.2300810, 0.3472850, 0.6168220, 0.4373380, 0.4581610, 0.9268800, 0.9311290, 0.7767140, 0.9376330, 0.6426660, 0.0735107, 0.1515400, 0.0839557, 0.1101690, 0.8279970, 0.9475250, 0.7580990, 0.4197480, 0.5121400, 0.9318340, 0.9723980, 0.0488850, 0.1443600, 0.8329140, 0.6298940, 0.7773880, 0.7867590, 0.5620150, 0.9461870, 0.0963216, 0.5817330, 0.5228370, 0.2059600, 0.6081160, 0.2050000, 0.4948940, 0.0860958, 0.1286550, 0.6540260, 0.9815180, 0.2869970, 0.7358540, 0.1517190, 0.4603600, 0.9076880, 0.8408280, 0.7902430, 0.6066630, 0.6041770, 0.2616000, 0.2493380, 0.9681610, 0.0243756, 0.1683480, 0.6549440, 0.3146720, 0.8983130, 0.2785320, 0.1638970, 0.3041480, 0.8968040, 0.2474500, 0.8736040, 0.9217050, 0.2073240, 0.1581440, 0.8274000, 0.8175310, 0.0209652, 0.6170280, 0.7712340, 0.2463910, 0.4992430, 0.6485610, 0.6824840, 0.0662828, 0.5006270, 0.5901800, 0.8065790, 0.1619750, 0.8923560, 0.8989150, 0.3405810, 0.3665800, 0.6583360, 0.8773270, 0.3062590, 0.2840300, 0.5034220, 0.7553370, 0.2520040, 0.7838800, 0.6576320, 0.5924670, 0.2518220, 0.0222373, 0.9754700, 0.4792720, 0.5831800, 0.3127430, 0.9505580, 0.7636070, 0.0740627, 0.8203380, 0.6932600, 0.8473530, 0.4511260, 0.7325800, 0.8695080, 0.4294500, 0.8497300, 0.0244342, 0.7438890, 0.1153210, 0.5367110, 0.5594470, 0.6417490, 0.4656020, 0.5371170, 0.5442880, 0.9679960, 0.8696190, 0.6447200, 0.9710580, 0.4860230, 0.0981751, 0.5203980, 0.4944520, 0.0287237, 0.3591480, 0.3448280, 0.3949690, 0.4683380, 0.9271290, 0.4746430, 0.5503100, 0.6845250, 0.3100160, 0.5004860, 0.3085530, 0.5125660, 0.5172720, 0.5782930, 0.7395950, 0.7401120, 0.2011690, 0.1888660, 0.7646220, 0.9406010, 0.7671510, 0.6974590, 0.4658760, 0.1449760, 0.0651553, 0.4508320, 0.9049640, 0.1573450, 0.7889830, 0.9666090, 0.9304070, 0.3273050, 0.3908870, 0.4926400, 0.6864060, 0.3740850, 0.8427110, 0.7769520, 0.2975730, 0.2836720, 0.1410290, 0.0471298, 0.2650680, 0.8761530, 0.1178040, 0.6045820, 0.0854878, 0.7922620, 0.9841660, 0.4793220, 0.4531850, 0.1551670, 0.9988600, 0.8598530, 0.0680528, 0.7690570, 0.6500170, 0.1105230, 0.5675370, 0.8412160, 0.5282070, 0.2260060, 0.7494560, 0.9775540, 0.6766340, 0.2892640, 0.4784970, 0.3278740, 0.6123010, 0.2511240, 0.5870870, 0.8185390, 0.5507540, 0.0649072, 0.6759200, 0.4078440, 0.6583410, 0.6082100, 0.1887670, 0.4723250, 0.3171130, 0.7999450, 0.8216430, 0.3717290, 0.5667140, 0.9183780, 0.3731090, 0.7516250, 0.2755580, 0.8547570, 0.8110810, 0.9542490, 0.5001440, 0.3627450, 0.3724250, 0.8639490, 0.8082350, 0.8683740, 0.6344900, 0.9433970, 0.7500870, 0.4346730, 0.2402820, 0.5409710, 0.1104140, 0.3150230, 0.6133970, 0.0429250, 0.6554340, 0.0769191, 0.5452300, 0.3200300, 0.4416860, 0.9030420, 0.4151380, 0.1384800, 0.6922410, 0.5702130, 0.5316730, 0.7473940, 0.3050970, 0.3390270, 0.2249470, 0.4946260, 0.1572370, 0.3329090, 0.2377060, 0.9026400, 0.3747280, 0.6090820, 0.3561800, 0.6995810, 0.0887090, 0.4660800, 0.0297640, 0.5890550, 0.3653020, 0.8800820, 0.3008230, 0.8009870, 0.1318400, 0.1841810, 0.2788460, 0.1089930, 0.1627880, 0.9749930, 0.7037380, 0.3012720, 0.3007340, 0.6580600, 0.9334450, 0.3836350, 0.6850360, 0.1118470, 0.0572202, 0.2049740, 0.8007940, 0.7879730, 0.5193340, 0.8869340, 0.9273160, 0.3099590, 0.3982700, 0.6612700, 0.4582260, 0.7986090, 0.6950680, 0.8233400, 0.5651030, 0.4829410, 0.6094470, 0.3298930, 0.4457500, 0.0581935, 0.7062700, 0.9848010, 0.9619890, 0.2694640, 0.4154770, 0.0733317, 0.6962590, 0.8005700, 0.8129610, 0.6659010, 0.4052400, 0.1568610, 0.6395730, 0.6897210, 0.5533670, 0.0755091, 0.9137180, 0.8709970, 0.3457780, 0.0523580, 0.0536171, 0.3302210, 0.9599850, 0.2757150, 0.8948740, 0.3899600, 0.8174190, 0.7841400, 0.7802590, 0.7058720, 0.4543660, 0.5034490, 0.3690840, 0.6152800, 0.8881320, 0.3071390, 0.5291240, 0.7426320, 0.8540270, 0.6004870, 0.3697830, 0.4892810, 0.8839950, 0.8280760, 0.7386410, 0.2745480, 0.7596200, 0.3244380, 0.1220780, 0.9236760, 0.4067570, 0.6527330, 0.1466220, 0.1196240, 0.8660100, 0.1989880, 0.8192890, 0.1952770, 0.9370270, 0.6238380, 0.0106947, 0.7564830, 0.8835870, 0.4755580, 0.4727840, 0.8561420, 0.1054790, 0.3820680, 0.2679930, 0.5900130, 0.9561380, 0.9572130, 0.1450420, 0.7136340, 0.7814420, 0.4969730, 0.5770190, 0.8577240, 0.9269110, 0.2646450, 0.1188250, 0.7516680, 0.8926410, 0.9175090, 0.3754880, 0.6493430, 0.4271670, 0.6204670, 0.3462960, 0.4498700, 0.2472510, 0.9473010, 0.6412720, 0.4701780, 0.5242390, 0.3242640, 0.1870650, 0.0697662, 0.3562780, 0.4601470, 0.9315170, 0.1895960, 0.0406114, 0.1927820, 0.0439304, 0.1135660, 0.7144200, 0.1179350, 0.8340060, 0.2107280, 0.2603290, 0.0726019, 0.4248550, 0.7532190, 0.3158730, 0.6141980, 0.2602430, 0.4236150, 0.0505977, 0.3829430, 0.5205280, 0.9537170, 0.0432796, 0.7368400, 0.2295840, 0.9270390, 0.3839860, 0.6024550, 0.2790830, 0.6796840, 0.6049910, 0.9279680, 0.1712960, 0.4532700, 0.6974550, 0.8082160, 0.0278487, 0.4382990, 0.0162567, 0.3509100, 0.5127270, 0.2382420, 0.5991990, 0.5369840, 0.9069510, 0.3706050, 0.2427140, 0.8264630, 0.1425730, 0.3464420, 0.9251850, 0.2422310, 0.5861260, 0.4973870, 0.1882990, 0.6603760, 0.7850910, 0.3268890, 0.4730780, 0.3508880, 0.7614440, 0.9258740, 0.1463590, 0.2942370, 0.0574084, 0.8680660, 0.2987980, 0.6423910, 0.0388906, 0.0488990, 0.0833396, 0.8873720, 0.1104880, 0.6413960, 0.4913440, 0.9128070, 0.4824740, 0.1130850, 0.1846420, 0.8097120, 0.8242290, 0.0804275, 0.0726569, 0.2693060, 0.9122380, 0.5440440, 0.9868730, 0.7465590, 0.6319780, 0.4040030, 0.7972480, 0.0242235, 0.2058630, 0.1962300, 0.6206010, 0.3998510, 0.6906880, 0.1840210, 0.1993480, 0.3358890, 0.3140590, 0.6742160, 0.0183406, 0.7248970, 0.6993930, 0.7935000, 0.7062070, 0.9834960, 0.9235670, 0.7301220, 0.7968760, 0.1971810, 0.5790670, 0.7999730, 0.0487226, 0.0819518, 0.0481986, 0.6664630, 0.9082780, 0.2515430, 0.4636100, 0.3983940, 0.1298460, 0.0031877, 0.4525190, 0.9113390, 0.8367810, 0.4966280, 0.8997650, 0.6329560, 0.6953330, 0.7260180, 0.2516330, 0.9697020, 0.5845420, 0.0958473, 0.4819440, 0.4616550, 0.7768150, 0.9534840, 0.4203930, 0.7242170, 0.2081550, 0.6274990, 0.3812210, 0.9641770, 0.6576710, 0.8011900, 0.7034320, 0.4219660, 0.0680710, 0.7285040, 0.3172720, 0.6674420, 0.8453970, 0.3938700, 0.1881790, 0.3771010, 0.0670405, 0.8355710, 0.8878290, 0.4031970, 0.0825356, 0.2749550, 0.7533860, 0.9710840, 0.3018420, 0.2917490, 0.1017570, 0.8530210, 0.2602370, 0.7335910, 0.7096800, 0.6860430, 0.0347647, 0.3806720, 0.6753870, 0.2315210, 0.2207330, 0.2122480, 0.6104220, 0.3803960, 0.6312920, 0.1610840, 0.3456540, 0.7016840, 0.8083950, 0.6746640, 0.2239380, 0.0883253, 0.8810600, 0.8147890, 0.2074880, 0.2852080, 0.6781970, 0.5960750, 0.3973330, 0.2559820, 0.5560350, 0.6168760, 0.2979160, 0.1689910, 0.6319160, 0.8960930, 0.2108200, 0.6992090, 0.0305803, 0.3650180, 0.1097590, 0.9313410, 0.0451927, 0.9432840, 0.7518910, 0.7120290, 0.4499930, 0.2604700, 0.7055650, 0.7867530, 0.6724280, 0.3155520, 0.9500930, 0.9771920, 0.9076350, 0.1692000, 0.1451780, 0.1513560, 0.7728630, 0.5820480, 0.9806020, 0.9672910, 0.9278470, 0.8619490, 0.2938910, 0.1427970, 0.6539070, 0.7886530, 0.8746680, 0.1799070, 0.7336360, 0.9921540, 0.1814080, 0.9732820, 0.1546490, 0.1371640, 0.9032230, 0.4512500, 0.7951920, 0.8124060, 0.6036310, 0.6600160, 0.2867620, 0.2232540, 0.7188420, 0.1479520, 0.0562004, 0.4389980, 0.3261980, 0.4921280, 0.9028780, 0.5741010, 0.7725160, 0.4437290, 0.6581610, 0.6564590, 0.7430420, 0.8951870, 0.9168820, 0.3124420, 0.4489630, 0.8235170, 0.3924410, 0.6673080, 0.4174260, 0.8154640, 0.3622960, 0.3895220, 0.5842470, 0.5729230, 0.5498000, 0.7444110, 0.8493200, 0.5539560, 0.7177360, 0.6562430, 0.8328810, 0.8589870, 0.4320050, 0.7794740, 0.8737130, 0.1860420, 0.7441080, 0.4379450, 0.4672380, 0.9781190, 0.3331110, 0.0069021, 0.6335920, 0.5756120, 0.7170400, 0.3932140, 0.2981410, 0.5433970, 0.7171390, 0.3388160, 0.8260560, 0.3419450, 0.0033949, 0.8800200, 0.3202740, 0.9717560, 0.2262490, 0.9917180, 0.2997350, 0.0725811, 0.0768797, 0.0171529, 0.0262706, 0.4371210, 0.1390850, 0.8516070, 0.5389780, 0.7017870, 0.1850610, 0.6852000, 0.7758230, 0.1757800, 0.7957140, 0.0267320, 0.8292540, 0.8756900, 0.8898390, 0.4484800, 0.8039610, 0.6930160, 0.3098020, 0.1123570, 0.8498750, 0.7541410, 0.6926730, 0.0667127, 0.7144230, 0.3379530, 0.1229840, 0.4772330, 0.8211490, 0.5217400, 0.8986580, 0.5373010, 0.9306720, 0.1246690, 0.9568210, 0.1993860, 0.5654370, 0.2575490, 0.5718070, 0.1258740, 0.3491750, 0.9668240, 0.2922710, 0.4113780, 0.1088470, 0.8790080, 0.4573400, 0.9124770, 0.3861000, 0.3834660, 0.1009920, 0.2578380, 0.3680490, 0.8026810, 0.4061390, 0.4868070, 0.3050680, 0.7831740, 0.5715400, 0.1442600, 0.0143831, 0.5403790, 0.6327030, 0.2130890, 0.1760800, 0.7957060, 0.9354280, 0.0982717, 0.6886910, 0.6059160, 0.4153910, 0.0161617, 0.9371400, 0.4902440, 0.9115290, 0.8039370, 0.5814260, 0.2819790, 0.4487670, 0.9555630, 0.4553150, 0.3252250, 0.2401600, 0.8837050, 0.2333170, 0.6790730, 0.9240630, 0.4622370, 0.9056040, 0.2065640, 0.9303700, 0.8063740, 0.2106900, 0.6936830, 0.0107263, 0.2704430, 0.8188470, 0.1254790, 0.6460690, 0.3639180, 0.0682959, 0.0879014, 0.7777810, 0.4056350, 0.4210820, 0.6780410, 0.5510330, 0.2701380, 0.9927700, 0.4328410, 0.1036720, 0.9590500, 0.2183040, 0.9714520, 0.7500960, 0.0886620, 0.4708780, 0.6583130, 0.0886299, 0.5299010, 0.1115630, 0.0549732, 0.4757100, 0.4442200, 0.2543620, 0.6448090, 0.2361610, 0.6098660, 0.4042710, 0.3309430, 0.0685391, 0.6891100, 0.9999000, 0.2608390, 0.9575180, 0.5937200, 0.2801520, 0.9472100, 0.9930840, 0.2698420, 0.5029350, 0.6442160, 0.6631220, 0.9944860, 0.1843600, 0.9026180, 0.3045040, 0.3770100, 0.0994732, 0.7317050, 0.2597950, 0.6499600, 0.7022950, 0.9681330, 0.7267770, 0.1524850, 0.1425540, 0.9156270, 0.7488130, 0.3994660, 0.0314711, 0.5459070, 0.5017350, 0.9943500, 0.7417070, 0.3910490, 0.2556370, 0.5187530, 0.4163890, 0.4187650, 0.1581000, 0.5196250, 0.6037380, 0.3598980, 0.8562940, 0.0754020, 0.5719880, 0.1851700, 0.1096140, 0.7150970, 0.4467230, 0.8067940, 0.2733800, 0.1537080, 0.2819410, 0.2649350, 0.1838230, 0.3200720, 0.7380300, 0.7429360, 0.6407590, 0.9951780, 0.2021160, 0.1433010, 0.4392840, 0.3941200, 0.0046220, 0.0410964, 0.0138828, 0.8597220, 0.9389250, 0.6629480, 0.8351270, 0.3983020, 0.1729690, 0.1551130, 0.7342880, 0.2129580, 0.0934144, 0.4835880, 0.2514890, 0.5794940, 0.7051220, 0.1659440, 0.0233259, 0.6631650, 0.3905510, 0.8030040, 0.1074270, 0.1628670, 0.1023020, 0.7862600, 0.3778650, 0.1177480, 0.7314530, 0.5506120, 0.9880990, 0.5601770, 0.8860170, 0.7258850, 0.4757080, 0.5371650, 0.2513310, 0.4604060, 0.5146120, 0.1061430, 0.8121900, 0.4632740, 0.8057070, 0.8913190, 0.9143180, 0.0765420, 0.9236730, 0.4701600, 0.4991830, 0.2504670, 0.4932760, 0.3200570, 0.3702420, 0.1238680, 0.6400160, 0.3038960, 0.8859340, 0.9783390, 0.7038970, 0.3754120, 0.5934700, 0.5454200, 0.9173110, 0.7968290, 0.2572130, 0.0170092, 0.8478990, 0.3311580, 0.1818790, 0.7147770, 0.3561890, 0.1113380, 0.9610210, 0.8832900, 0.1364800, 0.1031830, 0.1820840, 0.6006770, 0.7421890, 0.5808180, 0.9719610, 0.9820880, 0.7485840, 0.8235050, 0.8546100, 0.3614100, 0.4403330, 0.3039820, 0.2855840, 0.8044730, 0.7873650, 0.8227920, 0.0999929, 0.0107490, 0.6714590, 0.9013610, 0.2413730, 0.7020160, 0.9147280, 0.5269690, 0.7693590, 0.4322810, 0.1723690, 0.6909480, 0.6823750, 0.5152980, 0.1606530, 0.7041370, 0.2960450, 0.2794870, 0.3519860, 0.7324880, 0.3402170, 0.3637300, 0.2066360, 0.0088459, 0.9377250, 0.7604450, 0.9689850, 0.8851130, 0.4037620, 0.5513320, 0.3087420, 0.0410934, 0.2782170, 0.7897080, 0.2280890, 0.5199300, 0.5888680, 0.7933310, 0.4804210, 0.2747770, 0.6064480, 0.9957390, 0.2115140, 0.0714793, 0.1374840, 0.1902400, 0.8242220, 0.7209400, 0.1696830, 0.3515760, 0.8545110, 0.6802780, 0.4263660, 0.1247310, 0.9366150, 0.7823080, 0.5035770, 0.4191580, 0.3785110, 0.7005130, 0.8459220, 0.1965890, 0.8436730, 0.2465780, 0.0568229, 0.0886364, 0.9742390, 0.6604400, 0.1394270, 0.9525110, 0.0798754, 0.7465190, 0.3900440, 0.1101540, 0.6264880, 0.9260060, 0.0022569, 0.1985300, 0.0371682, 0.1820270, 0.4131950, 0.3779760, 0.7003410, 0.4439830, 0.2867850, 0.4439280, 0.6612380, 0.0739466, 0.2356560, 0.7328170, 0.4190720, 0.4270870, 0.4178020, 0.3349630, 0.7473100, 0.7366120, 0.1846120, 0.1511900, 0.6838920, 0.9722350, 0.3396160, 0.5906980, 0.2074520, 0.2579660, 0.4372480, 0.9735780, 0.7621780, 0.6030280, 0.7620650, 0.4071750, 0.6906480, 0.4385290, 0.3567640, 0.2972540, 0.1409800, 0.3846490, 0.4251900, 0.1895050, 0.2258070, 0.0964231, 0.7376100, 0.9657130, 0.4558040, 0.5428730, 0.2961420, 0.8113120, 0.4222870, 0.0521258, 0.8649540, 0.4469320, 0.6053590, 0.8683310, 0.8913260, 0.4156250, 0.7363210, 0.3184130, 0.9414810, 0.8948950, 0.0196171, 0.1934150, 0.3697680, 0.7886800, 0.6903130, 0.5380460, 0.1186170, 0.1799850, 0.4713690, 0.9215490, 0.5307660, 0.6789210, 0.7691720, 0.0448384, 0.0751929, 0.4623650, 0.7542800, 0.3210270, 0.6739340, 0.0953499, 0.2457920, 0.7227050, 0.7790460, 0.9969920, 0.0851839, 0.0515807, 0.7414000, 0.5814680, 0.6002550, 0.2489970, 0.0313345, 0.6589070, 0.6909210, 0.3687530, 0.0955238, 0.4568070, 0.2225270, 0.9636120, 0.2938860, 0.8580890, 0.0269452, 0.2233570, 0.7632270, 0.2244900, 0.7342310, 0.7131830, 0.6814350, 0.4452160, 0.0792896, 0.3053140, 0.3484530, 0.9336170, 0.1940700, 0.2674070, 0.9845280, 0.1990380, 0.5384300, 0.1418540, 0.2784150, 0.6316890, 0.8128160, 0.3014310, 0.1417590, 0.4541330, 0.4599450, 0.7649700, 0.0608002, 0.5903040, 0.7656660, 0.5711480, 0.2813780, 0.6662660, 0.6065650, 0.8585450, 0.5319080, 0.5840610, 0.9851040, 0.3061630, 0.5972500, 0.0577663, 0.1637810, 0.0154772, 0.0659443, 0.9380200, 0.2408390, 0.7813030, 0.7431930, 0.4463890, 0.0371092, 0.2966830, 0.3367490, 0.7797820, 0.7986120, 0.4617040, 0.4595280, 0.6891770, 0.5468210, 0.0304364, 0.4574750, 0.5820390, 0.1265660, 0.5027890, 0.2413280, 0.8223420, 0.1458870, 0.0650080, 0.3589850, 0.4959470, 0.4460890, 0.9570570, 0.4122600, 0.2733160, 0.7086590, 0.4812120, 0.8482060, 0.0836540, 0.3864750, 0.0572112, 0.4454990, 0.9290880, 0.9934440, 0.0559935, 0.4848310, 0.5453640, 0.6580150, 0.4052400, 0.7256200, 0.6117290, 0.5528620, 0.1966990, 0.4320750, 0.3105010, 0.2375020, 0.9673390, 0.0418932, 0.4324760, 0.9262060, 0.2570060, 0.1752810, 0.2884750, 0.9327030, 0.7207160, 0.1839590, 0.3390290, 0.0355379, 0.2472530, 0.1338200, 0.3517630, 0.4372010, 0.7347570, 0.5991290, 0.5575860, 0.6232130, 0.9048440, 0.4366180, 0.0673538, 0.4238680, 0.3712380, 0.6735120, 0.8677510, 0.5996860, 0.6005860, 0.8316980, 0.6517100, 0.2356120, 0.1331080, 0.6569190, 0.9444140, 0.3046250, 0.7248070, 0.6938310, 0.1341060, 0.1784080, 0.8263390, 0.8845620, 0.1157980, 0.0085163, 0.0901216, 0.6806320, 0.0894926, 0.6143570, 0.9543230, 0.4208310, 0.4759840, 0.2221050, 0.3163060, 0.5916320, 0.6003850, 0.5128670, 0.6036790, 0.3155650, 0.8554180, 0.2748680, 0.5939320, 0.2642890, 0.7253320, 0.8884430, 0.7861380, 0.7690330, 0.4821720, 0.8774940, 0.7783690, 0.8727020, 0.4709700, 0.6624940, 0.5645170, 0.3605270, 0.0209843, 0.0238200, 0.7764840, 0.3606660, 0.6537330, 0.5725100, 0.9205590, 0.8774330, 0.2377660, 0.3232430, 0.6927500, 0.8995140, 0.8502030, 0.3851060, 0.1449670, 0.7805980, 0.7653000, 0.0441152, 0.9460220, 0.6267420, 0.0401100, 0.8661000, 0.4472760, 0.9485800, 0.4144320, 0.8353030, 0.3843050, 0.4329110, 0.5086400, 0.3971780, 0.2517060, 0.9144290, 0.7624090, 0.1866000, 0.5076510, 0.3034740, 0.7416820, 0.3483210, 0.8965370, 0.8980950, 0.3382190, 0.9248320, 0.4188760, 0.9670120, 0.3581070, 0.2611760, 0.5183190, 0.8836680, 0.5033160, 0.7655010, 0.1468120, 0.7606490, 0.2072890, 0.6762170, 0.0041827, 0.6587590, 0.4470300, 0.0019818, 0.2026050, 0.5397070, 0.8762670, 0.2319790, 0.3918630, 0.8372900, 0.5978920, 0.1657670, 0.1834900, 0.9572890, 0.2477190, 0.9159290, 0.9027690, 0.3147300, 0.5140220, 0.3518530, 0.0200426, 0.7780180, 0.9472160, 0.6999110, 0.2189340, 0.0341567, 0.2463630, 0.7025040, 0.8532150, 0.7688320, 0.5697480, 0.5643410, 0.9587370, 0.2961780, 0.6975790, 0.4308970, 0.9274740, 0.2017700, 0.1076110, 0.8713550, 0.5393810, 0.1652670, 0.2738630, 0.4078490, 0.9192530, 0.5275350, 0.9298270, 0.1881680, 0.9036660, 0.9108320, 0.8730650, 0.5314270, 0.0762005, 0.1957790, 0.7385370, 0.9984160, 0.9432790, 0.4326940, 0.2475610, 0.4494540, 0.3918230, 0.0765929, 0.5121150, 0.4644510, 0.8389810, 0.8852800, 0.4374630, 0.0259770, 0.9487850, 0.6052520, 0.5603220, 0.6427070, 0.8134470, 0.1100770, 0.0404665, 0.5021050, 0.2044900, 0.5704570, 0.6502140, 0.6743960, 0.5259560, 0.9083330, 0.5319150, 0.2292480, 0.9499480, 0.3205930, 0.1610610, 0.7587440, 0.1691630, 0.0774608, 0.9042010, 0.0630772, 0.4468080, 0.9657350, 0.7953080, 0.4950440, 0.3146700, 0.7347300, 0.7311320, 0.9235100, 0.3088160, 0.1813920, 0.7017410, 0.3380940, 0.4399060, 0.2266030, 0.0192432, 0.6027730, 0.0299396, 0.5000990, 0.6345200, 0.4981350, 0.6117710, 0.4705240, 0.9121360, 0.3526160, 0.4861940, 0.5986130, 0.8167630, 0.6851240, 0.3576430, 0.7404680, 0.0993856, 0.8249710, 0.5559720, 0.6310030, 0.5496580, 0.7502190, 0.8236630, 0.1125720, 0.4738000, 0.7194930, 0.7162700, 0.8615780, 0.9304580, 0.1728590, 0.3050320, 0.6350060, 0.9821620, 0.9387950, 0.9640550, 0.9085050, 0.5922030, 0.7096800, 0.0641187, 0.2350920, 0.4631730, 0.1314030, 0.3308470, 0.3452190, 0.3849470, 0.9104590, 0.5117480, 0.9039060, 0.7834510, 0.9409220, 0.9154700, 0.1185240, 0.9024590, 0.1942500, 0.8772550, 0.8256450, 0.0264315, 0.9687750, 0.1044300, 0.5010490, 0.9860190, 0.3405150, 0.9012640, 0.2393320, 0.0418835, 0.5679730, 0.3448290, 0.9309690, 0.4839670, 0.3098120, 0.2463210, 0.2863000, 0.2770020, 0.4109560, 0.7062980, 0.2460370, 0.5948550, 0.1762920, 0.4067140, 0.8542300, 0.3955750, 0.5881530, 0.1540070, 0.7446510, 0.6260260, 0.7407620, 0.2242280, 0.2354440, 0.1773710, 0.2932310, 0.3993630, 0.9848360, 0.7853060, 0.0715314, 0.4583470, 0.1475050, 0.3539420, 0.6269660, 0.4942810, 0.8786880, 0.1518980, 0.1759810, 0.6040470, 0.2948180, 0.0221139, 0.3405480, 0.9505010, 0.1249950, 0.2343660, 0.8311120, 0.7880150, 0.4273130, 0.1519710, 0.6661210, 0.6168940, 0.9356340, 0.3398140, 0.7635060, 0.7552210, 0.7192920, 0.5066210, 0.8084800, 0.7013330, 0.7201260, 0.3998460, 0.2998730, 0.2121810, 0.6726600, 0.3253960, 0.8907460, 0.8964960, 0.3826920, 0.9223310, 0.9151190, 0.9307370, 0.4045500, 0.0303245, 0.7076940, 0.9208990, 0.9442710, 0.1036240, 0.4628940, 0.9155400, 0.4713100, 0.0586333, 0.0501928, 0.6003030, 0.1697000, 0.8249810, 0.1628220, 0.3120960, 0.5596870, 0.0998627, 0.9537050, 0.0670984, 0.2606090, 0.8015930, 0.4958000, 0.2081060, 0.3757080, 0.0465951, 0.8471300, 0.5806360, 0.4109030, 0.1774460, 0.6626860, 0.2796350, 0.5647750, 0.9155030, 0.0054472, 0.1353300, 0.9646300, 0.6092940, 0.1983000, 0.2614900, 0.3437160, 0.5179290, 0.5330650, 0.1488960, 0.3601810, 0.1859800, 0.1479270, 0.5967410, 0.1641880, 0.0077439, 0.1084440, 0.7409090, 0.1521720, 0.6397730, 0.2166450, 0.2528770, 0.5787550, 0.2044770, 0.2409870, 0.5726580, 0.1129180, 0.0904415, 0.6275460, 0.2796530, 0.5434550, 0.0544811, 0.1188550, 0.0460330, 0.3748390, 0.2871960, 0.9659730, 0.2169650, 0.0451074, 0.9725390, 0.3384610, 0.8002910, 0.4365440, 0.2841980, 0.7128300, 0.4725720, 0.5140350, 0.6957510, 0.2665670, 0.1873160, 0.5591180, 0.4419200, 0.2533530, 0.8203460, 0.9834950, 0.4049270, 0.0682481, 0.4201320, 0.6090930, 0.8750500, 0.5368220, 0.0651647, 0.0884921, 0.5782770, 0.9564990, 0.0962949, 0.3976800, 0.9778950, 0.7804310, 0.7718340, 0.9625710, 0.8331400, 0.6414430, 0.1591910, 0.9789260, 0.5816990, 0.5955090, 0.6397000, 0.6696080, 0.8337360, 0.5155240, 0.2084940, 0.1728470, 0.9008030, 0.7611310, 0.0175034, 0.4865220, 0.8029200, 0.5591900, 0.2937680, 0.3043240, 0.6629580, 0.2485120, 0.0089851, 0.2678110, 0.6410440, 0.6071410, 0.1430380, 0.9940510, 0.6165240, 0.8004630, 0.8732800, 0.2070050, 0.9197200, 0.4832290, 0.1799070, 0.8176040, 0.4347270, 0.3934950, 0.6269570, 0.9450710, 0.1962750, 0.8979280, 0.5453940, 0.4300720, 0.2847610, 0.4977820, 0.4143120, 0.6949330, 0.5262730, 0.6550410, 0.2456240, 0.0720961, 0.0672525, 0.1230230, 0.7243660, 0.8826410, 0.1079130, 0.3405130, 0.2291110, 0.1464050, 0.9819480, 0.0131648, 0.3813230, 0.5230450, 0.1936820, 0.6839650, 0.2358890, 0.8161990, 0.3079240, 0.0485912, 0.9768770, 0.4913760, 0.7979890, 0.8267090, 0.1977320, 0.0966480, 0.5245390, 0.9568630, 0.9487210, 0.0320569, 0.4941450, 0.9249160, 0.0236679, 0.5330130, 0.4324540, 0.0199176, 0.1281940, 0.5871840, 0.9718100, 0.2427310, 0.0173210, 0.5683740, 0.8913760, 0.9345810, 0.9108930, 0.8892280, 0.0120050, 0.2869960, 0.5677370, 0.7285800, 0.3474690, 0.0248862, 0.8164190, 0.5940750, 0.1143660, 0.4985940, 0.2020520, 0.0101962, 0.0811175, 0.7737780, 0.3058850, 0.1854430, 0.3821970, 0.2609950, 0.1327780, 0.6299630, 0.5734990, 0.2711470, 0.8297650, 0.1645060, 0.1034110, 0.9050790, 0.9609330, 0.5897560, 0.5237290, 0.1442120, 0.9769140, 0.4564110, 0.6168770, 0.3937040, 0.6681390, 0.6134640, 0.9176650, 0.9707330, 0.9287660, 0.7332660, 0.0520994, 0.0971854, 0.6078390, 0.6639340, 0.7251920, 0.9829830, 0.3577580, 0.3951110, 0.7950130, 0.1257370, 0.9097830, 0.0086155, 0.4026040, 0.1001930, 0.1620990, 0.0626661, 0.2889990, 0.3713030, 0.9231190, 0.9759580, 0.0184144, 0.3716330, 0.3127360, 0.9726110, 0.3837940, 0.1466290, 0.6576420, 0.8473160, 0.2984400, 0.2240340, 0.9330720, 0.0923674, 0.1391240, 0.4033710, 0.6058700, 0.9937500, 0.5639900, 0.0353394, 0.7769780, 0.4463610, 0.5038250, 0.3325170, 0.4872040, 0.6475260, 0.8071850, 0.7991180, 0.1048170, 0.2122110, 0.4261480, 0.2047180, 0.1125440, 0.6902530, 0.6519350, 0.2097800, 0.8649170, 0.5930900, 0.3528810, 0.3322690, 0.7775450, 0.3674470, 0.8020850, 0.5295660, 0.9575930, 0.0290406, 0.3045940, 0.8340010, 0.4451400, 0.7368430, 0.0838125, 0.2894720, 0.2658990, 0.8554380, 0.6793370, 0.0137773, 0.5798850, 0.4824830, 0.1509350, 0.1434640, 0.6789340, 0.7822420, 0.0369014, 0.4478720, 0.9979370, 0.2099570, 0.5928520, 0.6650950, 0.0832508, 0.9970340, 0.8002820, 0.9776120, 0.9649470, 0.8023790, 0.2137390, 0.3001240, 0.7580630, 0.1245510, 0.8326220, 0.7121580, 0.0580663, 0.0255578, 0.7956880, 0.8645920, 0.6069150, 0.1454470, 0.7286390, 0.4740050, 0.9489630, 0.4326320, 0.1530900, 0.2509080, 0.5831880, 0.6612920, 0.5570420, 0.5238200, 0.8987820, 0.2221830, 0.2003360, 0.0593240, 0.9263930, 0.1102600, 0.3897020, 0.1675870, 0.8639140, 0.3614660, 0.2368060, 0.2846520, 0.6749200, 0.3271200, 0.7953500, 0.0581647, 0.3651860, 0.7626500, 0.4797200, 0.0152387, 0.5184670, 0.5785580, 0.3152390, 0.7442630, 0.9479190, 0.1151660, 0.8151210, 0.9662070, 0.5899890, 0.6640540, 0.0293857, 0.5396030, 0.9215540, 0.3752010, 0.3628040, 0.7130540, 0.5606290, 0.1143230, 0.3620990, 0.6625100, 0.6960930, 0.3195310, 0.4907980, 0.6447710, 0.3864750, 0.4192400, 0.4434190, 0.8347110, 0.5943740, 0.4997970, 0.4770790, 0.3026320, 0.2937040, 0.7335020, 0.5039540, 0.2655760, 0.1436410, 0.3826160, 0.1556100, 0.9472350, 0.1354090, 0.1247010, 0.8675110, 0.3661300, 0.9542080, 0.1792590, 0.8244700, 0.7245860, 0.1617230, 0.6292700, 0.3263390, 0.9426320, 0.1088030, 0.6994210, 0.5134940, 0.7947810, 0.6203760, 0.2195040, 0.1287930, 0.8025950, 0.5741980, 0.6619960, 0.5545070, 0.8243980, 0.3858550, 0.0033573, 0.0879514, 0.6624150, 0.6435650, 0.8850400, 0.7254430, 0.9540330, 0.3923820, 0.3971860, 0.9080330, 0.3103020, 0.5761890, 0.0719431, 0.5836660, 0.5386110, 0.0319477, 0.2335920, 0.8674470, 0.3191750, 0.3448240, 0.1751720, 0.4685190, 0.8876720, 0.4213790, 0.4145860, 0.8573140, 0.4323740, 0.3765240, 0.0097540, 0.8255310, 0.4992480, 0.4555720, 0.3794920, 0.5479230, 0.4638370, 0.3782290, 0.8517690, 0.9340350, 0.7828310, 0.7179000, 0.0064826, 0.5836210, 0.0020279, 0.6691820, 0.0150271, 0.8437810, 0.6572440, 0.3472390, 0.2296570, 0.3900040, 0.2830420, 0.5064790, 0.2927160, 0.3231630, 0.6286390, 0.2051550, 0.0625641, 0.3572090, 0.2931580, 0.6233660, 0.9130940, 0.6137910, 0.6891480, 0.7996700, 0.6727560, 0.0740717, 0.0161664, 0.2382830, 0.4894200, 0.6345670, 0.8616890, 0.3743410, 0.8685630, 0.0868568, 0.2528890, 0.3467390, 0.6680280, 0.2316800, 0.3585670, 0.0070456, 0.5415430, 0.2845800, 0.4474190, 0.0161277, 0.6179950, 0.8977780, 0.8267580, 0.7684670, 0.0673586, 0.7255180, 0.2627280, 0.1800250, 0.0693277, 0.3949200, 0.0276382, 0.7401360, 0.2587430, 0.8778290, 0.1591590, 0.0590079, 0.6682420, 0.8249630, 0.4750070, 0.0953993, 0.2908360, 0.9944650, 0.5227340, 0.2103520, 0.0543161, 0.8273610, 0.8559850, 0.8714640, 0.5787530, 0.0739971, 0.3528260, 0.9101870, 0.3691620, 0.8005090, 0.3831430, 0.1487680, 0.7098080, 0.1718850, 0.4824220, 0.6074170, 0.0900390, 0.9905600, 0.5952870, 0.8006000, 0.3387680, 0.8800730, 0.0668824, 0.0619793, 0.2458950, 0.6719930, 0.1301810, 0.3508590, 0.7666160, 0.2812550, 0.5283090, 0.1853910, 0.4936180, 0.1404210, 0.1657940, 0.1615850, 0.2425020, 0.2677840, 0.4391080, 0.2171500, 0.2045150, 0.7062680, 0.4671380, 0.1701550, 0.1972820, 0.1029470, 0.9921230, 0.5983500, 0.1208110, 0.6812080, 0.2516800, 0.5865790, 0.7588460, 0.2641260, 0.0687151, 0.8161100, 0.1685730, 0.8792190, 0.9965600, 0.5815330, 0.4192180, 0.5710560, 0.0373040, 0.6226800, 0.2462770, 0.9228610, 0.8213840, 0.8353710, 0.7189620, 0.8265200, 0.6334370, 0.7047600, 0.3284800, 0.0992508, 0.9999430, 0.5281760, 0.2580850, 0.8896290, 0.4216660, 0.2180550, 0.4654220, 0.7291890, 0.3445350, 0.0410281, 0.4741960, 0.6940600, 0.5443700, 0.4999310, 0.2720250, 0.8194630, 0.2841660, 0.2053770, 0.2233730, 0.5304720, 0.8154390, 0.4137610, 0.7855550, 0.6149560, 0.3487740, 0.1968110, 0.6027300, 0.5156830, 0.2877520, 0.9323830, 0.3047330, 0.1329230, 0.4296720, 0.0791398, 0.5181630, 0.6290650, 0.5741080, 0.0445228, 0.4141000, 0.3401030, 0.8251790, 0.1156480, 0.4503550, 0.0384935, 0.2650700, 0.6768210, 0.3954580, 0.6340860, 0.8108140, 0.4910710, 0.6824350, 0.0527371, 0.9058190, 0.8097310, 0.2936430, 0.1323420, 0.0060620, 0.2155320, 0.3929310, 0.8689760, 0.2078710, 0.5470900, 0.9188020, 0.8952500, 0.0238992, 0.9070630, 0.8837090, 0.4138000, 0.2804270, 0.3386520, 0.9847680, 0.5867920, 0.4224510, 0.2607410, 0.1772300, 0.4791300, 0.5468170, 0.1584240, 0.9180220, 0.2061080, 0.8514860, 0.3706560, 0.2428500, 0.8482810, 0.6424020, 0.1859640, 0.2543820, 0.5797100, 0.5616820, 0.8238470, 0.4425880, 0.5871860, 0.1983230, 0.2108210, 0.4434370, 0.6174480, 0.9048640, 0.5833100, 0.6457910, 0.2527470, 0.2498470, 0.3442990, 0.0307163, 0.1198120, 0.5265200, 0.3213380, 0.1120410, 0.4543840, 0.4412560, 0.2518340, 0.1542250, 0.8838200, 0.1504580, 0.1868760, 0.9023180, 0.1693090, 0.6481940, 0.5582790, 0.2012620, 0.4743270, 0.1042210, 0.0192794, 0.9948370, 0.1753810, 0.7206320, 0.3256090, 0.6158460, 0.2121730, 0.2932340, 0.2288790, 0.8484120, 0.8931550, 0.1265640, 0.3602780, 0.1329450, 0.0961252, 0.4531660, 0.9460350, 0.6737610, 0.3587220, 0.5785800, 0.6340420, 0.2671750, 0.1317970, 0.0795050, 0.4006430, 0.9004260, 0.8722740, 0.5287980, 0.2602220, 0.8174870, 0.3065700, 0.0161465, 0.8567930, 0.4541920, 0.8394220, 0.7324600, 0.9832780, 0.4928540, 0.3007590, 0.7516540, 0.5821790, 0.5854110, 0.3560190, 0.5393120, 0.1436270, 0.4862220, 0.1761440, 0.4665770, 0.0461700, 0.3314950, 0.7618110, 0.9854230, 0.6386400, 0.8145440, 0.6714030, 0.6051770, 0.4260080, 0.9626790, 0.3561900, 0.8207280, 0.8369160, 0.9061150, 0.3617890, 0.2171260, 0.7065620, 0.8340940, 0.6537760, 0.6159830, 0.3738710, 0.9428040, 0.1093250, 0.3853150, 0.9932020, 0.2266780, 0.5011430, 0.3232160, 0.5303540, 0.8649110, 0.7433500, 0.1682300, 0.6432580, 0.9254050, 0.1762280, 0.6820240, 0.6198520, 0.0343160, 0.0219379, 0.0403421, 0.2438860, 0.8334350, 0.3595740, 0.9314520, 0.1431300, 0.2369550, 0.1889440, 0.9377620, 0.6214750, 0.0256183, 0.1703710, 0.0059248, 0.9546900, 0.3663640, 0.6809820, 0.2464190, 0.9386140, 0.0450350, 0.1778620, 0.0826315, 0.5820020, 0.6917680, 0.7232230, 0.6738070, 0.3630290, 0.5503760, 0.2320910, 0.2731440, 0.3324290, 0.3796900, 0.0500004, 0.2600680, 0.8270780, 0.8878490, 0.9999380, 0.3653450, 0.6736740, 0.2659990, 0.0257342, 0.7970330, 0.0190322, 0.6042010, 0.1973500, 0.9717630, 0.4098170, 0.2212930, 0.8752470, 0.9893220, 0.8366800, 0.7624480, 0.1372310, 0.0471065, 0.2562090, 0.6775220, 0.4292480, 0.5987920, 0.0364445, 0.0546215, 0.1505900, 0.2694830, 0.9335770, 0.8410180, 0.7991540, 0.0463197, 0.7172210, 0.8428970, 0.8876610, 0.5471570, 0.7654010, 0.3240370, 0.6042520, 0.6522300, 0.5221350, 0.3994190, 0.6210830, 0.4476930, 0.2534960, 0.6049630, 0.0992850, 0.6278080, 0.7117320, 0.3984240, 0.7731050, 0.5390240, 0.5791240, 0.7042540, 0.0537839, 0.6395220, 0.9673020, 0.9516410, 0.1149410, 0.7379500, 0.2336460, 0.8349190, 0.4822560, 0.9123790, 0.8875120, 0.2618580, 0.3185510, 0.9193270, 0.6465670, 0.3712800, 0.9338120, 0.8515290, 0.7182030, 0.0633297, 0.2104410, 0.6271090, 0.3453400, 0.8607250, 0.7858080, 0.8450850, 0.0757396, 0.4226110, 0.5353670, 0.1034970, 0.3818890, 0.5087040, 0.0982833, 0.5008450, 0.1614410, 0.8987060, 0.4922040, 0.7185780, 0.7575900, 0.3785120, 0.8798620, 0.6272630, 0.0859322, 0.0831147, 0.7199020, 0.1470350, 0.8801670, 0.2158210, 0.9451090, 0.3559600, 0.3943170, 0.4469060, 0.7815100, 0.3493570, 0.2484780, 0.6765630, 0.6506030, 0.0165982, 0.8380560, 0.6384810, 0.8257160, 0.6508040, 0.2253290, 0.0091007, 0.7248970, 0.2083120, 0.5803110, 0.0363395, 0.5160860, 0.2541450, 0.3582950, 0.4181650, 0.6330780, 0.1896670, 0.4610870, 0.1831760, 0.1414690, 0.5267000, 0.9532090, 0.6451680, 0.7629850, 0.6628050, 0.2988190, 0.8326820, 0.8669020, 0.0938690, 0.7075920, 0.4029380, 0.9954380, 0.0354619, 0.1219210, 0.8509270, 0.0205986, 0.3934930, 0.6015500, 0.0283034, 0.0681924, 0.9721320, 0.9663500, 0.9129590, 0.0801279, 0.9703010, 0.0740595, 0.5435100, 0.0413437, 0.2284550, 0.2616930, 0.2593970, 0.9337720, 0.1818030, 0.3176120, 0.9851080, 0.6060320, 0.8646740, 0.0600194, 0.8084490, 0.3806570, 0.4378470, 0.7311040, 0.2619230, 0.3102100, 0.6710820, 0.3459340, 0.1248930, 0.7235100, 0.4507480, 0.2863880, 0.3848510, 0.2076880, 0.1054770, 0.0408976, 0.8230150, 0.4289400, 0.4818640, 0.3026260, 0.8631110, 0.8262770, 0.6311690, 0.9935190, 0.5613400, 0.5059400, 0.0760910, 0.5325930, 0.0528393, 0.8390820, 0.4904090, 0.7447540, 0.3444270, 0.3853160, 0.3023220, 0.8964600, 0.1560410, 0.0019387, 0.8420880, 0.5270720, 0.6511450, 0.9936500, 0.2051980, 0.1472720, 0.4554400, 0.9045250, 0.4972440, 0.1200630, 0.8014430, 0.1509540, 0.2866620, 0.3030020, 0.1506150, 0.5002620, 0.8490060, 0.1048700, 0.4278870, 0.6358970, 0.5729400, 0.6033300, 0.6248430, 0.5842180, 0.9322160, 0.6684160, 0.8559760, 0.1087170, 0.1391850, 0.6603640, 0.8503390, 0.1158060, 0.0471439, 0.6862480, 0.8945030, 0.0557540, 0.1239850, 0.5289650, 0.9649080, 0.4059290, 0.1154080, 0.7772430, 0.0705450, 0.4534570, 0.0424666, 0.4129890, 0.5927890, 0.7860130, 0.2193540, 0.6525760, 0.4797930, 0.3651930, 0.0785947, 0.3982370, 0.7819590, 0.2818350, 0.4451710, 0.7657940, 0.4439270, 0.8982090, 0.8678350, 0.6211370, 0.6564280, 0.3088140, 0.1572150, 0.0640174, 0.4083960, 0.1852530, 0.0163881, 0.8161480, 0.8763490, 0.8626010, 0.8069290, 0.5035710, 0.5358500, 0.1054130, 0.9208540, 0.9966060, 0.5434210, 0.0943357, 0.2454370, 0.8997510, 0.3320010, 0.7298300, 0.5173140, 0.0893856, 0.9432110, 0.9255760, 0.7907540, 0.9230040, 0.3257940, 0.8439820, 0.3486980, 0.0846243, 0.1046720, 0.1789440, 0.3372710, 0.0212000, 0.6199980, 0.7724620, 0.8763160, 0.3898170, 0.4941530, 0.0025634, 0.0864728, 0.0887194, 0.7477110, 0.3943740, 0.9481560, 0.0358106, 0.6420540, 0.5864840, 0.2463680, 0.6027470, 0.3281930, 0.6949800, 0.0455525, 0.3804770, 0.7159700, 0.7115530, 0.7393450, 0.3685900, 0.4863020, 0.8511710, 0.3363810, 0.5483970, 0.8609030, 0.1949330, 0.5305030, 0.9163350, 0.6265140, 0.2591980, 0.2547390, 0.5269070, 0.8835680, 0.5934880, 0.4948940, 0.1872600, 0.6306080, 0.5501960, 0.6202870, 0.4935090, 0.1904530, 0.6351530, 0.9388780, 0.8800480, 0.6202510, 0.9894420, 0.8661110, 0.0943328, 0.0447234, 0.5272760, 0.0172759, 0.2834570, 0.7871990, 0.5939460, 0.8414870, 0.6235360, 0.6413100, 0.7953460, 0.9455220, 0.9524180, 0.0398149, 0.4072140, 0.6200430, 0.4078100, 0.1081440, 0.4456660, 0.5940820, 0.3145220, 0.9738180, 0.9265030, 0.6942130, 0.7773880, 0.1125610, 0.0515372, 0.5347760, 0.2548590, 0.8314090, 0.4883810, 0.1358340, 0.0017803, 0.3419840, 0.6487210, 0.6151240, 0.5784370, 0.6387380, 0.3669510, 0.6066370, 0.4714840, 0.6691680, 0.5644440, 0.1073290, 0.9411840, 0.3319690, 0.8706400, 0.0429139, 0.7841500, 0.4006100, 0.7327240, 0.0628692, 0.9334200, 0.7613380, 0.4791090, 0.3831120, 0.8783970, 0.9479390, 0.5371510, 0.0309643, 0.7676850, 0.0978479, 0.8881380, 0.8346920, 0.7069580, 0.1825530, 0.0297133, 0.1711960, 0.4783070, 0.9184450, 0.5942600, 0.5661500, 0.1727450, 0.5566970, 0.4834540, 0.2899620, 0.3498700, 0.1613520, 0.9099270, 0.9025690, 0.3004010, 0.0096054, 0.3640300, 0.1135410, 0.0603813, 0.6505990, 0.6984290, 0.0742893, 0.4281570, 0.7988700, 0.6279260, 0.1119010, 0.7644520, 0.8893260, 0.7283190, 0.8385430, 0.8288530, 0.6276820, 0.8982790, 0.0399592, 0.4452350, 0.9583940, 0.0198001, 0.5606050, 0.0206969, 0.2451750, 0.9797650, 0.2791310, 0.4660250, 0.2316180, 0.6428400, 0.6252120, 0.8246030, 0.6802390, 0.7779040, 0.5675930, 0.9545740, 0.7933950, 0.4650080, 0.3419620, 0.1055720, 0.7309790, 0.4598160, 0.1294830, 0.9904350, 0.7221130, 0.8330500, 0.7637750, 0.6034630, 0.8755690, 0.0100109, 0.0440273, 0.4037010, 0.5584490, 0.9358830, 0.4206580, 0.9393280, 0.3049790, 0.4582100, 0.1605070, 0.8999390, 0.4679120, 0.0214801, 0.6068120, 0.8862330, 0.0346405, 0.3798650, 0.2546220, 0.2184360, 0.9184660, 0.4238780, 0.5650570, 0.9976990, 0.0066047, 0.2328760, 0.4395790, 0.9015000, 0.2444710, 0.7098630, 0.6598330, 0.3141400, 0.9054720, 0.1478990, 0.7557370, 0.7745350, 0.1500950, 0.3422510, 0.2333450, 0.8347080, 0.2096140, 0.2663740, 0.6894370, 0.7885040, 0.0349016, 0.1011140, 0.3559100, 0.3601710, 0.8109900, 0.7871510, 0.9104290, 0.8214570, 0.5472840, 0.0144379, 0.5618930, 0.2400610, 0.3726400, 0.1769010, 0.5854440, 0.2360770, 0.0995898, 0.4430790, 0.6989230, 0.6632480, 0.8584300, 0.4488510, 0.9770270, 0.8719010, 0.4309460, 0.0241010, 0.4137440, 0.4890580, 0.9590390, 0.1557520, 0.2280030, 0.8892650, 0.2861100, 0.7205980, 0.5403670, 0.1686760, 0.9486990, 0.2338550, 0.8678260, 0.7771080, 0.9117490, 0.9960810, 0.3873020, 0.6148890, 0.1176510, 0.9769270, 0.5707490, 0.8595370, 0.2537440, 0.4874530, 0.2209590, 0.8313050, 0.7883570, 0.4161540, 0.7802810, 0.4111470, 0.5308590, 0.3210660, 0.1849560, 0.2700060, 0.4303020, 0.9831890, 0.8089830, 0.3051350, 0.9424950, 0.7772830, 0.9955700, 0.7461960, 0.0917753, 0.9504580, 0.6871510, 0.1232670, 0.0778065, 0.2639000, 0.8206220, 0.8382570, 0.5132520, 0.5083110, 0.6025400, 0.9777860, 0.3042760, 0.5829670, 0.4160840, 0.1325400, 0.5709420, 0.0648527, 0.1572940, 0.9616650, 0.8916720, 0.7671700, 0.1385080, 0.5587350, 0.9291270, 0.8318470, 0.5303540, 0.4664690, 0.9472730, 0.8369260, 0.6391960, 0.9821400, 0.3579170, 0.7609330, 0.1824070, 0.5429590, 0.8920430, 0.0714057, 0.3250850, 0.4214250, 0.1910300, 0.1362490, 0.4235600, 0.7174050, 0.4290600, 0.4274910, 0.3510510, 0.2435920, 0.5117700, 0.0724274, 0.8972660, 0.1581910, 0.2957020, 0.8607110, 0.8472540, 0.3222920, 0.8962660, 0.1707720, 0.7649590, 0.6621990, 0.8461260, 0.5472760, 0.5781620, 0.3801360, 0.1290290, 0.7079000, 0.9889540, 0.9831780, 0.4614990, 0.9795520, 0.4260890, 0.4715760, 0.3154860, 0.3172130, 0.6337530, 0.6141150, 0.9370460, 0.6601590, 0.0814412, 0.8143570, 0.8800030, 0.6928500, 0.6602660, 0.6247250, 0.8172480, 0.9559740, 0.4020650, 0.8491980, 0.6875060, 0.2229250, 0.0322573, 0.6222410, 0.7696740, 0.9330540, 0.5358250, 0.2829230, 0.7111010, 0.3118820, 0.9479710, 0.1846930, 0.1050890, 0.3101840, 0.9307690, 0.0966038, 0.5496420, 0.0806931, 0.2547390, 0.8543130, 0.2683850, 0.7919370, 0.4373320, 0.4295160, 0.1284620, 0.4940330, 0.7388650, 0.5313260, 0.6595610, 0.0443600, 0.8948950, 0.2171210, 0.4397680, 0.9243470, 0.2935920, 0.4570980, 0.1889180, 0.4372020, 0.8827290, 0.3207860, 0.7651690, 0.7183120, 0.5867500, 0.5534180, 0.0937736, 0.5909840, 0.8658870, 0.7899070, 0.9430680, 0.1349300, 0.3269480, 0.9329180, 0.7229240, 0.9427980, 0.8107170, 0.5192590, 0.7913310, 0.9803990, 0.7701070, 0.2702340, 0.8088230, 0.2016110, 0.5796310, 0.8139560, 0.2215090, 0.1838000, 0.4455830, 0.1183150, 0.4740460, 0.7843940, 0.6162930, 0.1393880, 0.2194530, 0.2644580, 0.5718740, 0.1958440, 0.7193440, 0.2492980, 0.3324370, 0.3609700, 0.2121390, 0.1343050, 0.5492330, 0.6976540, 0.0617535, 0.7836080, 0.1502650, 0.5234820, 0.1476840, 0.7557570, 0.6545180, 0.2488260, 0.7539450, 0.3508110, 0.2051380, 0.5889180, 0.4218700, 0.3505790, 0.1877200, 0.8234210, 0.5177830, 0.4574400, 0.0463071, 0.0810333, 0.2318810, 0.7120620, 0.8087460, 0.9859780, 0.5282310, 0.5515430, 0.3690430, 0.6484360, 0.6378530, 0.5588120, 0.1622500, 0.4892150, 0.2203550, 0.9473750, 0.7778120, 0.6208610, 0.3583440, 0.2253810, 0.6215890, 0.9193390, 0.6559700, 0.3600850, 0.5561980, 0.8361350, 0.2561970, 0.2944350, 0.3864300, 0.3496890, 0.9144980, 0.6696810, 0.7588770, 0.3921980, 0.7787640, 0.3472750, 0.2312620, 0.4863940, 0.1751950, 0.8491340, 0.1586140, 0.5007670, 0.8083890, 0.4594220, 0.7187590, 0.7097420, 0.9838870, 0.8419030, 0.8249640, 0.6988880, 0.6204630, 0.6635640, 0.8539020, 0.6885600, 0.1450690, 0.4103480, 0.6600690, 0.6104840, 0.0069241, 0.1386380, 0.8712030, 0.3871160, 0.6760480, 0.4104540, 0.6524610, 0.9110710, 0.7105840, 0.7649720, 0.9010710, 0.5629410, 0.7918850, 0.3536460, 0.7282120, 0.3487240, 0.8175710, 0.4366210, 0.2337290, 0.4680480, 0.5651200, 0.1511810, 0.4325790, 0.8038340, 0.2343770, 0.4096660, 0.5341190, 0.5581050, 0.6450120, 0.8012760, 0.8192940, 0.3800940, 0.6738140, 0.4941190, 0.4533950, 0.6906670, 0.6901210, 0.2315310, 0.5015570, 0.1677710, 0.2763820, 0.2703020, 0.0682647, 0.2561160, 0.1658450, 0.7523900, 0.3054740, 0.6622890, 0.7973880, 0.9443070, 0.9104970, 0.9913830, 0.1451240, 0.4215220, 0.7808320, 0.8848130, 0.6513010, 0.8773470, 0.9042420, 0.1509240, 0.2417380, 0.3342060, 0.6196030, 0.5774500, 0.0876481, 0.8249990, 0.7285020, 0.9974510, 0.2812120, 0.1594120, 0.9467670, 0.2035710, 0.4318710, 0.8797180, 0.8050430, 0.3219850, 0.4868110, 0.2372860, 0.0242833, 0.3216230, 0.0230816, 0.9627910, 0.8685140, 0.3340940, 0.9091180, 0.0681088, 0.8488260, 0.2342080, 0.5812450, 0.0212128, 0.0167556, 0.0154778, 0.1483550, 0.2317310, 0.6523400, 0.9441910, 0.9129980, 0.2690970, 0.4437870, 0.4830820, 0.3451260, 0.3452420, 0.2973760, 0.5098450, 0.8130390, 0.7651390, 0.1596860, 0.2152950, 0.0554305, 0.5819630, 0.0642794, 0.4347550, 0.1351120, 0.7763480, 0.5868900, 0.6846040, 0.9135290, 0.9277870, 0.6589960, 0.7368230, 0.2481330, 0.5467030, 0.0058570, 0.4264310, 0.1009660, 0.7734650, 0.0775056, 0.0350232, 0.4232490, 0.1789420, 0.4299720, 0.1391750, 0.7106630, 0.0992646, 0.6439150, 0.8548020, 0.2694790, 0.2363700, 0.6844880, 0.7739030, 0.5165800, 0.8867670, 0.7932690, 0.7800150, 0.6978320, 0.7602880, 0.0974523, 0.5645120, 0.0120290, 0.1772220, 0.7201020, 0.5628110, 0.1115640, 0.0962819, 0.7060820, 0.9200400, 0.8597800, 0.3120860, 0.5063680, 0.1958670, 0.0736621, 0.2554720, 0.5875250, 0.5094770, 0.7238470, 0.5253150, 0.6639990, 0.8446450, 0.7707180, 0.4871590, 0.5046420, 0.7403330, 0.1224590, 0.0862872, 0.4580870, 0.1176220, 0.0764084, 0.1152150, 0.4000370, 0.5758960, 0.7287530, 0.8938260, 0.2338620, 0.5689030, 0.5745510, 0.7781440, 0.4860590, 0.0245012, 0.8520750, 0.7849700, 0.2359560, 0.8708340, 0.9877980, 0.7639760, 0.7347480, 0.9205750, 0.5405010, 0.9023610, 0.7061020, 0.9347110, 0.4358190, 0.8116780, 0.3235760, 0.8785870, 0.4480520, 0.5510860, 0.4363020, 0.4445560, 0.0390137, 0.2154890, 0.3633380, 0.0932000, 0.8301650, 0.2273040, 0.9569050, 0.6971870, 0.8327620, 0.2566980, 0.7022790, 0.6882910, 0.6922130, 0.0084350, 0.8168230, 0.1873930, 0.6373410, 0.4266560, 0.3358540, 0.4680280, 0.1274550, 0.5063150, 0.2970270, 0.4138010, 0.7315430, 0.3581830, 0.4243770, 0.2915290, 0.9772880, 0.2494720, 0.9321720, 0.1996230, 0.4636030, 0.5243910, 0.0821644, 0.7167800, 0.9960420, 0.9288060, 0.2729010, 0.4118590, 0.7703070, 0.7221640, 0.1289110, 0.1867200, 0.8009420, 0.2183760, 0.1265140, 0.7245950, 0.1533230, 0.6423080, 0.0602161, 0.2334890, 0.7720080, 0.6811740, 0.6233330, 0.0549233, 0.1301650, 0.7850700, 0.7133270, 0.9385290, 0.0434140, 0.4660120, 0.8961920, 0.1480730, 0.5573810, 0.3087680, 0.8073890, 0.7573800, 0.4041140, 0.3068880, 0.6195100, 0.2066660, 0.4734010, 0.6678540, 0.5834130, 0.3022440, 0.8070340, 0.7466360, 0.1593760, 0.3168670, 0.9036420, 0.8216830, 0.0088289, 0.1615140, 0.4865870, 0.1792180, 0.0221330, 0.1969800, 0.8150890, 0.9676600, 0.4646200, 0.7351320, 0.1381710, 0.8078010, 0.6703600, 0.3763120, 0.5821910, 0.7780600, 0.4667230, 0.1880800, 0.9447150, 0.5817660, 0.3193660, 0.8224020, 0.6203770, 0.7702110, 0.1234560, 0.4370070, 0.2719860, 0.4959270, 0.3779970, 0.7437970, 0.3121900, 0.8948620, 0.2661300, 0.1418210, 0.4816740, 0.4745270, 0.3748320, 0.5278980, 0.1997220, 0.0258984, 0.5394100, 0.3068690, 0.7201190, 0.9924930, 0.9385230, 0.0538650, 0.8108000, 0.4794400, 0.2614240, 0.5037450, 0.5044760, 0.7807460, 0.6989360, 0.2029770, 0.1091900, 0.8698820, 0.8452620, 0.6872610, 0.0338568, 0.3670240, 0.1912400, 0.6499030, 0.8463920, 0.9214460, 0.4920640, 0.3684740, 0.4080950, 0.8256590, 0.4091020, 0.8680570, 0.8460580, 0.1763750, 0.9698890, 0.1631320, 0.4694270, 0.7518540, 0.9056100, 0.8298270, 0.5371890, 0.7874390, 0.2255200, 0.3187470, 0.0564143, 0.3182760, 0.3571440, 0.2723940, 0.1149780, 0.2763030, 0.6598050, 0.7610610, 0.7969380, 0.2416750, 0.6381310, 0.8669820, 0.9460510, 0.3548410, 0.8396410, 0.9360880, 0.9373330, 0.7877280, 0.4167200, 0.0100310, 0.9777320, 0.0563947, 0.8327910, 0.3383720, 0.2479120, 0.9494310, 0.1837850, 0.6916730, 0.3508010, 0.7488960, 0.8654520, 0.7552270, 0.7530320, 0.8393290, 0.7355700, 0.7345290, 0.1221360, 0.5456470, 0.5322040, 0.0618523, 0.6168420, 0.2581390, 0.6070860, 0.2042230, 0.1616800, 0.3981640, 0.1791680, 0.0694356, 0.4154780, 0.5826090, 0.1770780, 0.8302080, 0.1239950, 0.7482460, 0.4115380, 0.7817180, 0.1428700, 0.0120378, 0.6501160, 0.9965590, 0.4753140, 0.8864510, 0.0737092, 0.0487168, 0.0889213, 0.2481570, 0.9958760, 0.3373930, 0.2906870, 0.8495930, 0.9611340, 0.2466180, 0.3818900, 0.7281210, 0.0666338, 0.2088970, 0.0594443, 0.8031450, 0.3331850, 0.1903870, 0.6428290, 0.9536090, 0.4282880, 0.6792580, 0.9172630, 0.2174560, 0.0312667, 0.3701330, 0.7165940, 0.5390540, 0.6792390, 0.1915930, 0.8880860, 0.0228037, 0.7551580, 0.7633760, 0.2529530, 0.2278990, 0.2630020, 0.4656570, 0.4996190, 0.5541990, 0.4328610, 0.9976520, 0.6655150, 0.1390140, 0.0489010, 0.8187190, 0.9189420, 0.7948870, 0.4140500, 0.2076350, 0.2134430, 0.6290680, 0.3278670, 0.7467500, 0.2460240, 0.7160860, 0.4312450, 0.8688980, 0.3302980, 0.8523970, 0.7543290, 0.3024710, 0.4111610, 0.1815080, 0.0696232, 0.5158990, 0.7614100, 0.6104040, 0.0443505, 0.7194470, 0.4853960, 0.1176130, 0.0398136, 0.7143920, 0.6039330, 0.5281820, 0.7844940, 0.2162110, 0.4479920, 0.5558240, 0.7789990, 0.5379130, 0.6393910, 0.1131910, 0.0183018, 0.9325020, 0.6431840, 0.6195000, 0.6062350, 0.2371300, 0.4076920, 0.7571220, 0.3195750, 0.3898210, 0.3776000, 0.1207560, 0.7887450, 0.3129850, 0.0535412, 0.0872410, 0.7781940, 0.9499090, 0.1619540, 0.0631321, 0.2885850, 0.5135030, 0.4819710, 0.0990283, 0.8327370, 0.2882850, 0.4108460, 0.1891370, 0.6362750, 0.3595420, 0.1346990, 0.7213560, 0.7327950, 0.3515260, 0.2755080, 0.8505950, 0.6301360, 0.2509920, 0.4095950, 0.8619100, 0.7392700, 0.5053420, 0.5104620, 0.0332784, 0.9403200, 0.8258110, 0.9772770, 0.9935070, 0.1274330, 0.2659550, 0.0645554, 0.7652450, 0.9832480, 0.2760640, 0.2366000, 0.1992010, 0.1691330, 0.3534090, 0.3606880, 0.3583280, 0.4667810, 0.4516650, 0.9601620, 0.5316080, 0.7051450, 0.6029910, 0.1441980, 0.0428755, 0.8546260, 0.3342860, 0.8671980, 0.0963536, 0.3139370, 0.7021110, 0.6763910, 0.3080320, 0.8800900, 0.4163150, 0.6273810, 0.8830330, 0.7643390, 0.8947190, 0.3721400, 0.8913340, 0.5859810, 0.7416290, 0.6231810, 0.7081430, 0.8023780, 0.5149130, 0.1008200, 0.9034750, 0.0866791, 0.6475090, 0.8573820, 0.2287160, 0.9576110, 0.7612680, 0.3632650, 0.5785490, 0.1029350, 0.8170970, 0.0472543, 0.9512340, 0.2029860, 0.5788380, 0.9612100, 0.3579380, 0.9401490, 0.5825570, 0.1269300, 0.2819940, 0.1525630, 0.6837960, 0.0397417, 0.2058030, 0.1428800, 0.3068190, 0.8580840, 0.8067710, 0.4143250, 0.6696630, 0.4035320, 0.3617590, 0.9263210, 0.8366960, 0.9772730, 0.3057590, 0.4090280, 0.1207940, 0.3393340, 0.1147090, 0.4969030, 0.7562670, 0.1254870, 0.0603031, 0.4278440, 0.3805690, 0.5127440, 0.5233840, 0.3530480, 0.3369950, 0.6686030, 0.5819150, 0.0944701, 0.6826070, 0.4623700, 0.7746240, 0.2146930, 0.0747197, 0.3460950, 0.9852300, 0.6761780, 0.4779500, 0.5046250, 0.4850180, 0.9100250, 0.3880090, 0.1104310, 0.9019600, 0.2057870, 0.0680880, 0.5197650, 0.5093110, 0.5181040, 0.6017500, 0.2643520, 0.8366960, 0.6419650, 0.1928490, 0.2599040, 0.6738210, 0.1621790, 0.7427590, 0.3748850, 0.3344950, 0.2208470, 0.7189280, 0.3769090, 0.2461170, 0.1716260, 0.8223960, 0.7547470, 0.0309723, 0.6670790, 0.0950698, 0.2410960, 0.5854040, 0.1811550, 0.7838770, 0.8423740, 0.2065630, 0.6818180, 0.7736710, 0.2845860, 0.5452980, 0.1704190, 0.9069140, 0.8026770, 0.7612390, 0.8105770, 0.9022610, 0.8922820, 0.9876480, 0.0551125, 0.9909280, 0.2705860, 0.8133470, 0.0401272, 0.5321470, 0.6710550, 0.1641830, 0.3340720, 0.0085984, 0.3955870, 0.5694100, 0.2058280, 0.6231630, 0.9592520, 0.6692020, 0.3651480, 0.8063640, 0.2298790, 0.2729340, 0.1152350, 0.1675660, 0.8025020, 0.8549110, 0.0927040, 0.5566110, 0.1210790, 0.5879580, 0.6284830, 0.5622470, 0.7840730, 0.0156109, 0.9702150, 0.2971000, 0.7872590, 0.0900517, 0.6404830, 0.6450400, 0.2741590, 0.4755660, 0.3239330, 0.8911380, 0.8629010, 0.0717405, 0.3708390, 0.4614970, 0.1920510, 0.4837260, 0.3569600, 0.7311950, 0.3940240, 0.5357190, 0.4332040, 0.7009750, 0.1955840, 0.7088830, 0.9032870, 0.9488750, 0.4558430, 0.2714140, 0.8061660, 0.2071390, 0.7993400, 0.3566810, 0.6395160, 0.6527850, 0.0329423, 0.4876070, 0.1654860, 0.1414310, 0.3793680, 0.8412030, 0.4305740, 0.1053830, 0.2825470, 0.4815080, 0.8660860, 0.7744450, 0.5634050, 0.6047410, 0.3985170, 0.8435070, 0.5977030, 0.7962340, 0.7678090, 0.2927970, 0.0254912, 0.8009740, 0.4411330, 0.4552920, 0.0399669, 0.4473230, 0.9811830, 0.9838710, 0.9087810, 0.1142110, 0.5185810, 0.3566110, 0.3254510, 0.3512860, 0.0853675, 0.2484180, 0.6869920, 0.5724860, 0.3979020, 0.2080640, 0.7154390, 0.7514400, 0.9234770, 0.0003031, 0.6962600, 0.2087630, 0.4196360, 0.1755100, 0.8507920, 0.1869600, 0.1054950, 0.9724310, 0.8909110, 0.9229360, 0.2167160, 0.8696740, 0.1965600, 0.1416850, 0.9287280, 0.1434960, 0.3968730, 0.8227110, 0.5207580, 0.8640350, 0.4519300, 0.9246130, 0.3358760, 0.7821630, 0.9320160, 0.1017900, 0.9264290, 0.5264240, 0.4805420, 0.6809750, 0.5298240, 0.7351360, 0.1617300, 0.2288170, 0.3819390, 0.2155930, 0.5953450, 0.0610633, 0.1088130, 0.1133930, 0.6972800, 0.7001680, 0.6156020, 0.5754820, 0.3628710, 0.2060510, 0.8322060, 0.7401250, 0.7296780, 0.9628790, 0.9747230, 0.1820070, 0.3384920, 0.1296980, 0.7973630, 0.1154980, 0.3624730, 0.8799620, 0.1258180, 0.2581920, 0.3391280, 0.5669700, 0.1302200, 0.1554500, 0.7798280, 0.2868660, 0.8375270, 0.9123270, 0.3923480, 0.7245090, 0.9207330, 0.4817710, 0.4563670, 0.7312880, 0.3942350, 0.3160820, 0.2945310, 0.7049150, 0.6758510, 0.4377490, 0.9553310, 0.1848050, 0.8544810, 0.3148030, 0.0179629, 0.0096313, 0.9784190, 0.1869520, 0.5388030, 0.7004060, 0.3307290, 0.5171580, 0.2552090, 0.0874535, 0.4594690, 0.3083320, 0.3006730, 0.6372100, 0.7344350, 0.1542220, 0.7329770, 0.2747430, 0.0412590, 0.3699940, 0.4339700, 0.6696260, 0.5962440, 0.4590540, 0.0402685, 0.2279560, 0.5526180, 0.8543610, 0.7522570, 0.8033170, 0.0913645, 0.3526500, 0.7795990, 0.3287460, 0.6182860, 0.6602400, 0.0129809, 0.2045170, 0.9994220, 0.3400840, 0.9797840, 0.3013910, 0.5790020, 0.9993470, 0.0416820, 0.9099070, 0.9060480, 0.8783200, 0.5856240, 0.5854260, 0.7667870, 0.1591330, 0.5568800, 0.3977360, 0.1785590, 0.6844520, 0.5138890, 0.7864510, 0.2567350, 0.4084750, 0.6296960, 0.9299140, 0.8172530, 0.1040890, 0.9713060, 0.4658630, 0.3005230, 0.9088880, 0.2408610, 0.2555380, 0.7496200, 0.7083390, 0.9015960, 0.2088700, 0.0546467, 0.7995540, 0.5420430, 0.9404770, 0.8833890, 0.4086490, 0.6914240, 0.2292370, 0.2959610, 0.4796300, 0.7699810, 0.9058370, 0.3255430, 0.6700960, 0.0293111, 0.3015610, 0.3065480, 0.3524530, 0.5605500, 0.0749766, 0.8530460, 0.7307560, 0.9814780, 0.7895130, 0.6394980, 0.9169800, 0.7473280, 0.3277930, 0.3880350, 0.7849900, 0.2624410, 0.6967140, 0.4078490, 0.8573450, 0.7022980, 0.8995020, 0.7391700, 0.4718250, 0.4265580, 0.5692760, 0.7056820, 0.3196560, 0.3878980, 0.9034150, 0.2622770, 0.8553990, 0.5606660, 0.1994190, 0.9431540, 0.2843240, 0.2631460, 0.1175740, 0.6572160, 0.3981360, 0.3218690, 0.7399040, 0.1272890, 0.6836330, 0.0443592, 0.5049820, 0.1052530, 0.4752400, 0.3488790, 0.9458880, 0.1307740, 0.0800247, 0.8699250, 0.7088820, 0.5921340, 0.5735460, 0.7032990, 0.1049670, 0.6744880, 0.9932830, 0.9406240, 0.6618750, 0.6546180, 0.6945160, 0.4330580, 0.1064470, 0.3842790, 0.6346170, 0.4275290, 0.0471097, 0.0389134, 0.8739330, 0.5458760, 0.3936490, 0.5082370, 0.6765930, 0.5076200, 0.1613650, 0.0646274, 0.5042640, 0.1198460, 0.9910640, 0.8978360, 0.2090020, 0.6461470, 0.4518270, 0.8630970, 0.4147070, 0.8147480, 0.6465180, 0.4168560, 0.4882770, 0.8256050, 0.2587430, 0.8552430, 0.2128310, 0.8418950, 0.2283450, 0.8106110, 0.9660030, 0.3880220, 0.2684760, 0.5002540, 0.5656540, 0.5841980, 0.6837030, 0.8271040, 0.9864020, 0.7721380, 0.3181270, 0.6600300, 0.8212050, 0.2643760, 0.4333430, 0.3421140, 0.5685010, 0.6075040, 0.2877150, 0.2209690, 0.6928810, 0.8229160, 0.0686032, 0.4527980, 0.7500290, 0.6078230, 0.7196200, 0.7272130, 0.9937990, 0.0885869, 0.7160500, 0.3948080, 0.5152490, 0.7246290, 0.1149850, 0.8788800, 0.3282080, 0.4042060, 0.8055170, 0.2917970, 0.2770590, 0.3688060, 0.5688550, 0.0494264, 0.2521430, 0.5569780, 0.4678540, 0.2954490, 0.7406270, 0.7139830, 0.7006790, 0.7049090, 0.3780840, 0.3656010, 0.0377609, 0.2022980, 0.1862930, 0.8647790, 0.4868630, 0.1398640, 0.8318760, 0.5195110, 0.0417034, 0.1889850, 0.3834040, 0.2394200, 0.5430350, 0.0330618, 0.8404620, 0.1276510, 0.7758110, 0.2477380, 0.5804330, 0.1155220, 0.3322140, 0.0312512, 0.1078060, 0.2747860, 0.7611560, 0.6334190, 0.0792952, 0.2097830, 0.2619090, 0.1416330, 0.7249750, 0.0826577, 0.3259170, 0.2591940, 0.4837790, 0.2496080, 0.6468570, 0.7710460, 0.6955040, 0.2178100, 0.7861590, 0.7966600, 0.1653980, 0.0579180, 0.3965800, 0.2956520, 0.3180380, 0.6872120, 0.8583670, 0.0100248, 0.6590500, 0.3656150, 0.1044960, 0.8798790, 0.2965540, 0.4197170, 0.7629680, 0.4993950, 0.5668400, 0.8134680, 0.7044340, 0.9994760, 0.8587120, 0.6391310, 0.3391040, 0.6912390, 0.2554010, 0.9803460, 0.2703110, 0.3301820, 0.6157730, 0.8092000, 0.2592160, 0.3343900, 0.7692690, 0.2113210, 0.2943610, 0.3362210, 0.3984000, 0.5138410, 0.9851810, 0.1481880, 0.7975630, 0.0772372, 0.5378400, 0.7942580, 0.8903600, 0.3019130, 0.1968840, 0.3169650, 0.6118480, 0.7314610, 0.5211760, 0.4488720, 0.1867550, 0.9255430, 0.9355850, 0.8451530, 0.5986100, 0.8828990, 0.2030960, 0.8319130, 0.8676280, 0.5379560, 0.8066510, 0.9718460, 0.8124200, 0.1732510, 0.2293380, 0.5281510, 0.2454710, 0.3496020, 0.5333120, 0.1877210, 0.9421160, 0.5232340, 0.9404880, 0.2738880, 0.6376560, 0.2160190, 0.3703260, 0.3749530, 0.1199610, 0.9348460, 0.0766564, 0.6990140, 0.0504058, 0.9383700, 0.2030210, 0.9905360, 0.6198280, 0.1559450, 0.4065230, 0.5677030, 0.3176260, 0.5019330, 0.3985410, 0.6928710, 0.5326770, 0.8355310, 0.8367460, 0.5104820, 0.1264810, 0.4886530, 0.6862370, 0.6949400, 0.7436030, 0.5069020, 0.4209610, 0.7028760, 0.2679320, 0.9210850, 0.8193200, 0.8573050, 0.6231690, 0.3579190, 0.8385110, 0.8915650, 0.8441850, 0.5166510, 0.8610100, 0.6461740, 0.7128950, 0.9023290, 0.8857160, 0.0898873, 0.1498220, 0.4722950, 0.9761220, 0.2166790, 0.6637250, 0.9080230, 0.2560590, 0.7637680, 0.6306360, 0.7114940, 0.9029620, 0.6934270, 0.1648630, 0.4171470, 0.2678000, 0.1668550, 0.5487790, 0.9206170, 0.5849850, 0.6555030, 0.5799730, 0.9629840, 0.5726740, 0.1245790, 0.4078350, 0.3576130, 0.7356340, 0.9212810, 0.7189050, 0.2084740, 0.1179450, 0.3389810, 0.3846310, 0.5123830, 0.8863940, 0.7319620, 0.3634050, 0.6735440, 0.7757880, 0.5235610, 0.0551718, 0.3654190, 0.4839470, 0.8763640, 0.1913520, 0.8505230, 0.4669870, 0.0122764, 0.4835110, 0.4900600, 0.8918090, 0.5797090, 0.6604110, 0.2759680, 0.6470600, 0.4610120, 0.8365240, 0.8881730, 0.1525530, 0.5338820, 0.7308340, 0.8923280, 0.0689471, 0.9244750, 0.3977590, 0.6045800, 0.8380910, 0.6339330, 0.7804400, 0.5259840, 0.0743586, 0.9223830, 0.0304374, 0.2556810, 0.5937160, 0.1990260, 0.3357470, 0.3354940, 0.8553910, 0.1440970, 0.2188270, 0.7550370, 0.8546720, 0.6852890, 0.9196570, 0.3773830, 0.8013930, 0.5072740, 0.6831440, 0.1898590, 0.3526240, 0.5121430, 0.0023810, 0.2450540, 0.1869620, 0.0394044, 0.1395390, 0.7391430, 0.1329890, 0.3127320, 0.5059450, 0.4072840, 0.8501430, 0.2086080, 0.3921570, 0.9286030, 0.5144600, 0.8848670, 0.6923290, 0.8465120, 0.0510279, 0.4682520, 0.2399980, 0.4404380, 0.9076860, 0.4076630, 0.7309700, 0.1321490, 0.3123980, 0.2496820, 0.7761620, 0.4308470, 0.3273610, 0.5942540, 0.2563940, 0.9725210, 0.2343570, 0.4181250, 0.0367356, 0.0002581, 0.7590680, 0.8925390, 0.6873600, 0.0632103, 0.4882050, 0.2925360, 0.0209426, 0.0319664, 0.3022910, 0.7390970, 0.8633650, 0.7177540, 0.2277430, 0.4996580, 0.9342170, 0.2821030, 0.7099330, 0.0663115, 0.3164920, 0.7927500, 0.7168020, 0.2896290, 0.3109150, 0.3322970, 0.4958980, 0.3798560, 0.3071810, 0.3202810, 0.1237270, 0.7711460, 0.2639300, 0.0393609, 0.4416580, 0.7757530, 0.8018970, 0.2836030, 0.3562680, 0.2486120, 0.9222900, 0.9373850, 0.5066950, 0.7759640, 0.8856900, 0.3911200, 0.9492350, 0.5335490, 0.2601940, 0.0242934, 0.1105210, 0.8060760, 0.1345330, 0.2366360, 0.5883350, 0.5700960, 0.1949760, 0.3286470, 0.3535620, 0.0252438, 0.8693100, 0.1919360, 0.1841560, 0.5306730, 0.8395020, 0.1029860, 0.8515620, 0.0073128, 0.9379520, 0.6891200, 0.4652800, 0.3604530, 0.0943165, 0.2143790, 0.1283890, 0.4404190, 0.3215570, 0.1033640, 0.2567640, 0.1121800, 0.8060430, 0.1830400, 0.0300327, 0.7981150, 0.0876145, 0.6078250, 0.6515060, 0.7852200, 0.0003939, 0.8564330, 0.1988760, 0.3473050, 0.2526030, 0.8032090, 0.0525653, 0.1601290, 0.5687110, 0.2064280, 0.8024060, 0.5510010, 0.6322040, 0.3645730, 0.8756230, 0.2273680, 0.3178610, 0.1142270, 0.2632640, 0.6889540, 0.7364390, 0.8566200, 0.7578180, 0.0027823, 0.7659730, 0.8210810, 0.7372870, 0.5950600, 0.1856710, 0.5461930, 0.8583560, 0.3745460, 0.3258360, 0.2717450, 0.4746340, 0.5074710, 0.9854870, 0.7881150, 0.7590720, 0.5843330, 0.4396570, 0.5718110, 0.2361060, 0.5025100, 0.4605100, 0.5814340, 0.0266095, 0.2769300, 0.0600933, 0.8588990, 0.1549260, 0.9093580, 0.3860420, 0.6943550, 0.3205350, 0.4390410, 0.7775050, 0.8548950, 0.0438629, 0.9745560, 0.7586800, 0.0942665, 0.6994600, 0.6906070, 0.3436720, 0.7670220, 0.8642510, 0.3078370, 0.8471620, 0.6470330, 0.0384919, 0.0048546, 0.1297930, 0.6274050, 0.5444790, 0.4406800, 0.6645930, 0.1879670, 0.2700100, 0.1144110, 0.1744320, 0.3377750, 0.9331380, 0.1758950, 0.3250600, 0.8248690, 0.1173480, 0.6585420, 0.3743110, 0.1430970, 0.1727050, 0.4937330, 0.3224860, 0.1047000, 0.9496920, 0.8479470, 0.0733369, 0.4996690, 0.1515700, 0.2415230, 0.7386220, 0.9106520, 0.9409610, 0.0002451, 0.4118850, 0.2796310, 0.8343080, 0.9131970, 0.0712455, 0.7768410, 0.7548610, 0.7422630, 0.5729370, 0.2597440, 0.3280320, 0.2594420, 0.9826500, 0.5235960, 0.0630599, 0.0842793, 0.4208610, 0.1498110, 0.9945200, 0.0900374, 0.7260670, 0.2544050, 0.1778420, 0.8532840, 0.6555360, 0.8788600, 0.8166150, 0.3617300, 0.0844249, 0.1451790, 0.7310030, 0.3230100, 0.8652150, 0.1865830, 0.9537770, 0.7791130, 0.1011690, 0.5195360, 0.4074110, 0.1800210, 0.0111473, 0.9774200, 0.8708810, 0.5855090, 0.1383760, 0.8679270, 0.9992430, 0.4370080, 0.1688650, 0.6617430, 0.5923540, 0.8104060, 0.4780900, 0.8426090, 0.5154680, 0.4989420, 0.8991020, 0.8449300, 0.2248270, 0.9732260, 0.5115070, 0.8377550, 0.3958110, 0.3535680, 0.1704790, 0.0933160, 0.6268000, 0.4725360, 0.3512600, 0.3276800, 0.6651800, 0.9674340, 0.0759273, 0.9447610, 0.7506850, 0.1003290, 0.5099460, 0.6718810, 0.0782687, 0.5980920, 0.0763919, 0.9155680, 0.7790510, 0.5832020, 0.1096420, 0.7761810, 0.8892880, 0.6681260, 0.9729910, 0.4074770, 0.5251620, 0.6405740, 0.5398890, 0.7099540, 0.5999780, 0.7151920, 0.2943340, 0.0468385, 0.7610180, 0.0137457, 0.3893830, 0.8282940, 0.8756390, 0.4473690, 0.5946320, 0.9825290, 0.3523460, 0.6292290, 0.4474920, 0.7967050, 0.0143345, 0.2179750, 0.4333680, 0.7121570, 0.3097470, 0.2759670, 0.8319890, 0.2795420, 0.7756620, 0.8070530, 0.5804890, 0.5556610, 0.5962280, 0.7781850, 0.7627890, 0.2148710, 0.6262220, 0.8588200, 0.3804160, 0.1277000, 0.7780480, 0.0102694, 0.2740060, 0.7808250, 0.6460470, 0.8151640, 0.7114730, 0.8204370, 0.9073380, 0.4555840, 0.9566050, 0.2094050, 0.9197860, 0.3682960, 0.1540830, 0.6048200, 0.2726530, 0.9193520, 0.6524970, 0.8631760, 0.9527650, 0.2331530, 0.4174820, 0.9911360, 0.8587820, 0.2348230, 0.6245360, 0.4820730, 0.7667600, 0.0746647, 0.7099110, 0.6322260, 0.9344820, 0.2986130, 0.3561330, 0.5688840, 0.4491680, 0.7856750, 0.1311950, 0.4301250, 0.1397590, 0.3748160, 0.5064210, 0.6700600, 0.4219150, 0.0565923, 0.9240160, 0.7499240, 0.3853460, 0.3988590, 0.5466820, 0.5676310, 0.6860200, 0.3388120, 0.1520210, 0.8699250, 0.5501580, 0.0884858, 0.0707294, 0.0360947, 0.9925940, 0.1151390, 0.5430990, 0.4035510, 0.1653590, 0.9553290, 0.3128270, 0.7347880, 0.4463560, 0.3482750, 0.7947380, 0.7073550, 0.3597570, 0.4287990, 0.1333090, 0.0469885, 0.4946730, 0.6040520, 0.8060650, 0.8899190, 0.9576460, 0.5710340, 0.1123520, 0.7159980, 0.1207080, 0.7575870, 0.7153000, 0.5660780, 0.0741200, 0.9267540, 0.5097280, 0.9592180, 0.3126450, 0.1555260, 0.9516400, 0.6616650, 0.6547590, 0.3617900, 0.0913561, 0.6167760, 0.3131100, 0.0889531, 0.7091380, 0.8379560, 0.5838240, 0.7119300, 0.8088880, 0.0098490, 0.0442400, 0.1079240, 0.9960040, 0.6567110, 0.7250290, 0.5285420, 0.9144590, 0.1806840, 0.6256780, 0.6927580, 0.7114560, 0.5125150, 0.4942970, 0.1300690, 0.9398510, 0.7238170, 0.0539918, 0.1251040, 0.4064620, 0.2776410, 0.3290520, 0.4914960, 0.7041290, 0.4319360, 0.4018740, 0.2629730, 0.3444160, 0.7303450, 0.2039170, 0.8682480, 0.1143580, 0.9632970, 0.5723690, 0.1703170, 0.2210410, 0.4696560, 0.0367894, 0.4901100, 0.8438520, 0.0336523, 0.4349650, 0.5984840, 0.7361900, 0.4479080, 0.1468940, 0.0537699, 0.4361360, 0.9025110, 0.3317730, 0.4942650, 0.9049310, 0.5037500, 0.4612410, 0.0131670, 0.0796726, 0.1371710, 0.4772460, 0.5706540, 0.5569830, 0.2397630, 0.0681506, 0.7441910, 0.1965010, 0.4392790, 0.2475710, 0.2442170, 0.6872640, 0.8309630, 0.0943247, 0.6855990, 0.6314490, 0.6934840, 0.3156020, 0.6188160, 0.6504480, 0.7689640, 0.9759620, 0.9431210, 0.2734060, 0.6916870, 0.2829780, 0.7405780, 0.5132710, 0.2840720, 0.8466270, 0.4377440, 0.1293580, 0.8634750, 0.5181350, 0.4180970, 0.4672970, 0.6661440, 0.9307510, 0.9328480, 0.8434240, 0.2038370, 0.0484700, 0.0654234, 0.2435460, 0.5770140, 0.2272430, 0.6503990, 0.1457640, 0.7123330, 0.8461200, 0.0769397, 0.0027125, 0.1804890, 0.4721980, 0.0537011, 0.8307480, 0.6984510, 0.9185610, 0.1438220, 0.9462780, 0.5501270, 0.4344660, 0.8745370, 0.2432950, 0.2766450, 0.4190360, 0.5773160, 0.1695910, 0.5727230, 0.5385260, 0.8102600, 0.4765700, 0.6296730, 0.9466230, 0.0911797, 0.9582610, 0.3060180, 0.2489480, 0.2980160, 0.6543960, 0.7313460, 0.1908050, 0.6299890, 0.1314200, 0.6054080, 0.6553020, 0.0392747, 0.0016036, 0.8118200, 0.0439506, 0.2244210, 0.6246460, 0.2002010, 0.0604689, 0.6623970, 0.5894860, 0.7270430, 0.9483980, 0.7608160, 0.3625070, 0.9787240, 0.8167640, 0.0194039, 0.0363092, 0.9046650, 0.7696150, 0.1721170, 0.4299730, 0.0375507, 0.9591010, 0.4357310, 0.8256210, 0.7619370, 0.6559900, 0.8274090, 0.3075210, 0.7531700, 0.4386050, 0.1186800, 0.2164860, 0.8733930, 0.4350720, 0.5713110, 0.9589040, 0.1262940, 0.2126830, 0.0593809, 0.2970900, 0.5644690, 0.0661398, 0.5634560, 0.8244630, 0.0236241, 0.5926760, 0.5714910, 0.2210900, 0.7532510, 0.6757480, 0.6717270, 0.9466090, 0.3777130, 0.2180070, 0.9063860, 0.1212520, 0.1177930, 0.3833750, 0.3712170, 0.9562020, 0.1143080, 0.0625160, 0.8211020, 0.3745720, 0.8597470, 0.2654050, 0.0661358, 0.9070500, 0.2936510, 0.1448740, 0.6496710, 0.5760270, 0.1751090, 0.5556560, 0.5316600, 0.7871670, 0.4399240, 0.0495554, 0.2099670, 0.3059210, 0.2723860, 0.9469130, 0.8932170, 0.4011130, 0.2165730, 0.5789130, 0.8916140, 0.8794580, 0.6529360, 0.9849970, 0.9584060, 0.9665330, 0.6200810, 0.0852327, 0.8599370, 0.6510680, 0.0737527, 0.5256060, 0.4293400, 0.4898520, 0.0495969, 0.3316360, 0.1010360, 0.4305130, 0.4524610, 0.9970690, 0.9142950, 0.3897390, 0.1025270, 0.2709120, 0.9016920, 0.9284570, 0.7619350, 0.5004000, 0.8890190, 0.1740580, 0.4531650, 0.2751070, 0.5139180, 0.9094010, 0.1905540, 0.2484010, 0.1320920, 0.1651500, 0.9811360, 0.9333140, 0.2031540, 0.1247640, 0.9761730, 0.3753690, 0.7348820, 0.3186400, 0.9091480, 0.7446760, 0.4024290, 0.9333000, 0.5055510, 0.9073640, 0.8903580, 0.3033550, 0.6184700, 0.8678870, 0.8429220, 0.5121420, 0.0571880, 0.6495130, 0.0870660, 0.3602070, 0.1059940, 0.3323900, 0.5834250, 0.6011080, 0.6298900, 0.4705730, 0.5546600, 0.7899950, 0.4644170, 0.4847730, 0.9307950, 0.7098590, 0.3510430, 0.9279510, 0.9031290, 0.6913180, 0.8027630, 0.8104350, 0.0291575, 0.0424378, 0.9058840, 0.7367520, 0.7297060, 0.5716500, 0.5887730, 0.4524430, 0.7453440, 0.6724210, 0.6607100, 0.1292430, 0.2724230, 0.0583755, 0.2454840, 0.6804100, 0.6561430, 0.3566350, 0.5058380, 0.6771690, 0.2462740, 0.1714080, 0.3708150, 0.0307692, 0.9813320, 0.3672660, 0.8173590, 0.4568280, 0.8528000, 0.7633040, 0.6241410, 0.3205290, 0.0319117, 0.1397740, 0.0682755, 0.0593937, 0.1245380, 0.3881340, 0.4746570, 0.5340040, 0.6231320, 0.3757130, 0.8075130, 0.8319700, 0.8720440, 0.6383330, 0.1714290, 0.4989400, 0.7294840, 0.4260080, 0.4560860, 0.9122070, 0.3120810, 0.7215490, 0.8308060, 0.6361300, 0.2288080, 0.0049750, 0.3829750, 0.2530510, 0.3229160, 0.8982680, 0.2415750, 0.4703690, 0.9967360, 0.8801140, 0.4746960, 0.1786680, 0.4425230, 0.3202830, 0.8954500, 0.6990870, 0.3883720, 0.4944120, 0.5241670, 0.0916707, 0.6441680, 0.9987710, 0.7536180, 0.1485180, 0.9159330, 0.5575080, 0.0139027, 0.7817130, 0.9362350, 0.5090210, 0.8151030, 0.7432730, 0.0794652, 0.4551110, 0.5837320, 0.0209827, 0.9370470, 0.8664150, 0.6363650, 0.3051060, 0.9924930, 0.8166750, 0.5675280, 0.7221350, 0.5390160, 0.0834244, 0.7820070, 0.5421700, 0.6489020, 0.8037810, 0.3888970, 0.8281840, 0.9818040, 0.3863620, 0.8871410, 0.5191440, 0.1025780, 0.2004700, 0.3546830, 0.9454080, 0.4515680, 0.8602310, 0.0364347, 0.6787650, 0.9638370, 0.7753890, 0.1607060, 0.1319310, 0.9678830, 0.1231220, 0.3933760, 0.5865610, 0.0043871, 0.3478430, 0.8840700, 0.1982730, 0.6915600, 0.2884140, 0.3264780, 0.2157190, 0.4137260, 0.4398220, 0.5767100, 0.4160030, 0.3643500, 0.6541560, 0.3900680, 0.5853030, 0.2981270, 0.9264510, 0.3917510, 0.0672380, 0.1296370, 0.2519310, 0.0542657, 0.2104220, 0.7289580, 0.4465780, 0.8840550, 0.6598770, 0.9635920, 0.5902470, 0.4596630, 0.8628490, 0.2906810, 0.9853310, 0.4491930, 0.3812270, 0.9776520, 0.8578470, 0.3774990, 0.1314220, 0.3636730, 0.5341870, 0.6070450, 0.2885370, 0.1497940, 0.9590810, 0.3758630, 0.6867520, 0.6940700, 0.4970440, 0.4107060, 0.5279280, 0.1221210, 0.5027700, 0.0579641, 0.3515090, 0.6703620, 0.4365640, 0.1408700, 0.7758160, 0.6744640, 0.7426150, 0.9096980, 0.6183830, 0.1473980, 0.7721400, 0.2287250, 0.7642160, 0.6608350, 0.2455770, 0.3077000, 0.8999210, 0.2136990, 0.2722600, 0.5821470, 0.1121880, 0.6269650, 0.7701110, 0.4659950, 0.3989590, 0.0249761, 0.4608710, 0.7735710, 0.2882700, 0.4679220, 0.3986260, 0.2302170, 0.6828400, 0.9858600, 0.6744890, 0.7251850, 0.7659030, 0.5365550, 0.0388318, 0.2810960, 0.0094818, 0.1824000, 0.0543675, 0.4602130, 0.1594570, 0.1487300, 0.5671660, 0.5584570, 0.4901420, 0.4539740, 0.9551260, 0.0391636, 0.9147660, 0.5879850, 0.2210130, 0.6180760, 0.5591750, 0.1997880, 0.2411770, 0.2525980, 0.3595520, 0.7568810, 0.9911070, 0.8959230, 0.1680980, 0.4308860, 0.6261300, 0.4554410, 0.2206840, 0.4238250, 0.3449720, 0.5536400, 0.0834057, 0.0123263, 0.8786650, 0.5189500, 0.5947650, 0.4107980, 0.9470580, 0.5202570, 0.5844400, 0.5012810, 0.3560790, 0.1472540, 0.4792060, 0.2822230, 0.9387500, 0.6591090, 0.9694370, 0.3828870, 0.5535090, 0.7791630, 0.0060378, 0.7877350, 0.1822670, 0.0837992, 0.3869350, 0.4719070, 0.4729820, 0.6876510, 0.3976880, 0.1586570, 0.1474180, 0.3097190, 0.9066780, 0.5667820, 0.7388580, 0.1002350, 0.4825040, 0.9796110, 0.3585610, 0.6244030, 0.0673108, 0.3334340, 0.4548050, 0.8894740, 0.7910710, 0.5957500, 0.8371760, 0.6024830, 0.5636050, 0.3884330, 0.2622280, 0.8538550, 0.6585690, 0.8309260, 0.9159020, 0.2890140, 0.5671340, 0.3940770, 0.5744190, 0.4398010, 0.9688760, 0.2631710, 0.8821740, 0.0899146, 0.2423100, 0.1755870, 0.1473270, 0.3162260, 0.1345490, 0.4218410, 0.9575500, 0.9200490, 0.2217300, 0.0651255, 0.1898940, 0.1888670, 0.8752420, 0.1815470, 0.3103830, 0.6310760, 0.5129920, 0.5417190, 0.5246500, 0.7833460, 0.9709110, 0.5218430, 0.4237280, 0.5663710, 0.1560470, 0.3804560, 0.0795515, 0.1787340, 0.8199120, 0.9561220, 0.8601260, 0.7042560, 0.5986520, 0.5981860, 0.3251590, 0.8087790, 0.8859930, 0.1624810, 0.6396550, 0.5371420, 0.8041180, 0.6773600, 0.7105640, 0.9888750, 0.2421440, 0.1195680, 0.9901670, 0.8718140, 0.5734980, 0.9298440, 0.0768512, 0.6378220, 0.2196050, 0.6769110, 0.1198700, 0.5563150, 0.5194210, 0.6921240, 0.3123690, 0.2869880, 0.1926880, 0.5413320, 0.7083660, 0.4332520, 0.8095740, 0.5743500, 0.1918170, 0.9579990, 0.1428630, 0.5949110, 0.4371180, 0.3601980, 0.5379370, 0.0900658, 0.9806090, 0.2667910, 0.4626810, 0.6079800, 0.5483990, 0.3967000, 0.6605980, 0.9107110, 0.1618530, 0.6916620, 0.4194430, 0.9887750, 0.7095600, 0.5348310, 0.3829850, 0.5247720, 0.1942990, 0.0486218, 0.2346310, 0.4487720, 0.8875840, 0.9419500, 0.7061050, 0.8015130, 0.5049510, 0.7994130, 0.0993259, 0.4847890, 0.7608390, 0.7585490, 0.7503160, 0.6300580, 0.6077380, 0.0183900, 0.2036680, 0.0811137, 0.1620850, 0.5591340, 0.6648120, 0.4747380, 0.4965580, 0.2513120, 0.3586910, 0.8031020, 0.4020840, 0.1667460, 0.8114650, 0.6567600, 0.3818620, 0.6295030, 0.5949470, 0.9522160, 0.2152600, 0.3596580, 0.2096670, 0.0638479, 0.8524910, 0.6336740, 0.8762860, 0.9779700, 0.0717024, 0.3432200, 0.5815380, 0.3549950, 0.0240097, 0.3419940, 0.9567660, 0.9454150, 0.6839630, 0.4603400, 0.2054170, 0.2361750, 0.7881030, 0.3660830, 0.4813920, 0.0307963, 0.5668730, 0.9980950, 0.6760990, 0.5713710, 0.8709400, 0.2974750, 0.2519910, 0.6206930, 0.3328930, 0.3024220, 0.1227460, 0.3698760, 0.2366170, 0.3430080, 0.4252410, 0.8043420, 0.8502210, 0.5369490, 0.0731873, 0.3862450, 0.9580480, 0.4047870, 0.7634470, 0.1886960, 0.4104290, 0.2219820, 0.9891980, 0.2611010, 0.6515670, 0.3008280, 0.5792310, 0.1442000, 0.8713180, 0.0959588, 0.9092230, 0.8178780, 0.8938810, 0.1961980, 0.3286270, 0.7375050, 0.1463450, 0.3206360, 0.5252080, 0.8476610, 0.1264580, 0.1987050, 0.5917300, 0.7061830, 0.8712260, 0.0504174, 0.3625460, 0.3686920, 0.5678900, 0.3439400, 0.0266605, 0.8318670, 0.7030550, 0.7789620, 0.9877800, 0.3703470, 0.1448340, 0.5719560, 0.0314400, 0.9581170, 0.0367400, 0.7225930, 0.8519230, 0.3135890, 0.4274990, 0.3894370, 0.9665930, 0.5964330, 0.6087320, 0.0976957, 0.5371090, 0.2206840, 0.5741540, 0.3267780, 0.8207290, 0.8795720, 0.8802820, 0.6739120, 0.0792683, 0.7990430, 0.7078060, 0.6301340, 0.6496760, 0.4880430, 0.1980670, 0.7395490, 0.4464440, 0.1483460, 0.1011140, 0.3006310, 0.2661460, 0.7287140, 0.3517880, 0.5553930, 0.1496160, 0.6089140, 0.2596210, 0.5003860, 0.0087119, 0.9611300, 0.1340090, 0.7914530, 0.7333590, 0.2077890, 0.7513140, 0.0303066, 0.3291660, 0.9401660, 0.6132510, 0.7104850, 0.0873139, 0.0713638, 0.5251020, 0.9427210, 0.7539890, 0.2318640, 0.9508440, 0.0175312, 0.1753540, 0.7994040, 0.4428100, 0.4211750, 0.1339760, 0.3926920, 0.2449900, 0.5225230, 0.1474050, 0.9869860, 0.6657610, 0.2201630, 0.2396060, 0.9217890, 0.3316050, 0.3207950, 0.6727620, 0.8329010, 0.2681190, 0.2205900, 0.2070920, 0.4992470, 0.0783398, 0.0438265, 0.9931600, 0.5400090, 0.1067360, 0.7113940, 0.1640900, 0.2211650, 0.3030330, 0.6258770, 0.7620340, 0.9002250, 0.1555770, 0.0653495, 0.2855960, 0.7684040, 0.9864560, 0.6190280, 0.5045010, 0.0727039, 0.6965200, 0.4923440, 0.8624810, 0.5760120, 0.3837800, 0.2742440, 0.6007880, 0.9780910, 0.2981300, 0.4248160, 0.7105870, 0.6985420, 0.6542200, 0.6026190, 0.4233560, 0.2561030, 0.1764480, 0.5699280, 0.8558270, 0.3045680, 0.9287720, 0.8006500, 0.5894910, 0.8964780, 0.1094930, 0.7657240, 0.9452350, 0.1841590, 0.7682790, 0.7535330, 0.8518360, 0.4982770, 0.1536940, 0.3164090, 0.5424910, 0.7781440, 0.8832200, 0.1052730, 0.0789349, 0.5359890, 0.3270280, 0.1108620, 0.5597160, 0.0957215, 0.4685350, 0.5006760, 0.0561586, 0.4637200, 0.5447280, 0.9786200, 0.8275720, 0.3767410, 0.1337620, 0.6784660, 0.7782700, 0.5232390, 0.7042210, 0.5235920, 0.8727990, 0.4524660, 0.3249850, 0.0407172, 0.7428810, 0.5034350, 0.3944930, 0.3781150, 0.8895380, 0.2915700, 0.7752750, 0.3777380, 0.5162740, 0.5697020, 0.8168490, 0.2055100, 0.1596890, 0.3796380, 0.0049407, 0.2355350, 0.1936960, 0.2370800, 0.6929730, 0.7625020, 0.4736670, 0.6604500, 0.3896250, 0.2766280, 0.4455750, 0.9521720, 0.0438460, 0.8691520, 0.0886530, 0.5816130, 0.9248280, 0.8655590, 0.4137990, 0.3613810, 0.7354360, 0.0834471, 0.3772960, 0.6117360, 0.4750670, 0.9304720, 0.8958840, 0.9119970, 0.6443010, 0.7573790, 0.1751040, 0.4771960, 0.6075910, 0.0316759, 0.8909950, 0.7552540, 0.6013850, 0.4541480, 0.3001530, 0.1940150, 0.5679990, 0.3454210, 0.1206760, 0.4908340, 0.3517180, 0.6389950, 0.4865850, 0.9055510, 0.0349440, 0.7734500, 0.1027030, 0.8316530, 0.0476182, 0.7019470, 0.4668770, 0.5780800, 0.9716450, 0.7911880, 0.8202110, 0.0300508, 0.9304820, 0.8098760, 0.3722680, 0.1531660, 0.9140600, 0.1559740, 0.2092830, 0.8733940, 0.9439590, 0.2975400, 0.6088170, 0.7114110, 0.1130500, 0.6817640, 0.6717250, 0.5995870, 0.1593010, 0.4287520, 0.0608098, 0.7921680, 0.3166890, 0.0139623, 0.2030040, 0.6428640, 0.0959260, 0.8409980, 0.4153150, 0.5771820, 0.2536320, 0.4071960, 0.4041110, 0.7980820, 0.6626660, 0.6494940, 0.2812140, 0.5803290, 0.3979730, 0.3466190, 0.5256430, 0.7780970, 0.6962870, 0.9766260, 0.9878030, 0.7477770, 0.0231587, 0.9039560, 0.4688770, 0.1839870, 0.1844340, 0.1139650, 0.9600590, 0.5512250, 0.2032460, 0.6738480, 0.9428460, 0.1683600, 0.4660200, 0.7866360, 0.8060830, 0.8508210, 0.6104190, 0.4475630, 0.6624770, 0.8402560, 0.0367073, 0.0830511, 0.1882080, 0.3027520, 0.8022800, 0.4022110, 0.1412110, 0.5498220, 0.9796130, 0.9339470, 0.1928990, 0.9999170, 0.5494880, 0.6527960, 0.1788780, 0.1950270, 0.4725690, 0.4429590, 0.6442440, 0.7241710, 0.6857500, 0.3885870, 0.4842170, 0.4886960, 0.0959492, 0.8894800, 0.9443100, 0.8512380, 0.1264500, 0.0754582, 0.6067550, 0.0259175, 0.3880470, 0.0499229, 0.2315210, 0.5809180, 0.5933300, 0.9356580, 0.6238950, 0.9858270, 0.8320580, 0.4669860, 0.8792230, 0.9534090, 0.7899170, 0.9492450, 0.5929010, 0.7686030, 0.5298740, 0.3434300, 0.0020623, 0.8215180, 0.8906340, 0.5882500, 0.5869070, 0.6043460, 0.2353820, 0.3905920, 0.8506060, 0.8669460, 0.4985650, 0.4585210, 0.7070730, 0.7924890, 0.3385730, 0.8151940, 0.3160890, 0.5555250, 0.2921690, 0.7194840, 0.3252390, 0.6677750, 0.9800640, 0.8640280, 0.3971090, 0.1429820, 0.7707780, 0.1845100, 0.0672438, 0.9863180, 0.2005390, 0.4857420, 0.6208730, 0.3433090, 0.2244240, 0.4041550, 0.3522070, 0.0289449, 0.6930030, 0.1207300, 0.8441990, 0.5352490, 0.7087130, 0.8827450, 0.3514410, 0.3943530, 0.6366440, 0.7345230, 0.8476800, 0.8547430, 0.8652740, 0.9167470, 0.8462790, 0.7793750, 0.0216243, 0.5001630, 0.9640820, 0.9047080, 0.9337730, 0.7900020, 0.3816840, 0.6086670, 0.2442210, 0.6406890, 0.0591546, 0.0077804, 0.2844310, 0.3135140, 0.5112920, 0.0589001, 0.5612410, 0.9663400, 0.6476540, 0.4393670, 0.5162950, 0.6588760, 0.1004830, 0.7725110, 0.9611470, 0.9358730, 0.8601550, 0.2879840, 0.9316060, 0.7069210, 0.9802650, 0.9175620, 0.2690180, 0.7374460, 0.2463910, 0.3253590, 0.5922760, 0.3219660, 0.4443510, 0.6574920, 0.8857070, 0.9905100, 0.7750800, 0.8661510, 0.7186690, 0.3485740, 0.3469510, 0.8092120, 0.5228070, 0.7012910, 0.2332920, 0.8406170, 0.8420500, 0.0136862, 0.3779820, 0.7750910, 0.4492740, 0.4440760, 0.5588890, 0.8209210, 0.7129090, 0.5047320, 0.2656670, 0.0855162, 0.8893360, 0.2401450, 0.3738640, 0.0426084, 0.8631380, 0.8095200, 0.1679920, 0.4162240, 0.9089890, 0.8448830, 0.3432730, 0.7026890, 0.0327272, 0.1436760, 0.8260420, 0.7243670, 0.4331600, 0.9836830, 0.7473120, 0.7378360, 0.4397140, 0.0587682, 0.2654470, 0.4777810, 0.6739060, 0.7245950, 0.3549630, 0.3089220, 0.4911910, 0.3247700, 0.5402200, 0.4016140, 0.7269100, 0.2460220, 0.2400840, 0.3499660, 0.6175610, 0.4750530, 0.7838780, 0.5994620, 0.4724980, 0.6871560, 0.7768320, 0.7327190, 0.4510350, 0.1324150, 0.4858400, 0.4084630, 0.6163690, 0.0279878, 0.6692240, 0.2010270, 0.6217030, 0.0466045, 0.5903340, 0.1120810, 0.1115190, 0.6634830, 0.7596490, 0.7997920, 0.2345570, 0.7599040, 0.5265600, 0.2808400, 0.4959200, 0.4285870, 0.7677080, 0.2967350, 0.6234140, 0.6729430, 0.2890160, 0.9804940, 0.8630890, 0.4252500, 0.4544260, 0.1470540, 0.7182640, 0.7854770, 0.3644700, 0.1828140, 0.8038400, 0.3683900, 0.6843210, 0.7006640, 0.4368930, 0.9954650, 0.7993050, 0.3157050, 0.7084720, 0.7231870, 0.3601810, 0.5867270, 0.8597270, 0.0821735, 0.9423120, 0.6964310, 0.6871200, 0.2460860, 0.5722900, 0.0075383, 0.4780110, 0.2833940, 0.1681280, 0.7876420, 0.3360780, 0.4863470, 0.3976610, 0.0207008, 0.3549740, 0.6132670, 0.5116450, 0.3987060, 0.0850598, 0.6562250, 0.2778210, 0.2506990, 0.3523180, 0.0919646, 0.5613690, 0.4876360, 0.3054780, 0.6553880, 0.2869440, 0.2720080, 0.0048795, 0.1213200, 0.9582440, 0.3325230, 0.6453210, 0.3883660, 0.6052070, 0.9236080, 0.6565580, 0.3791070, 0.5542680, 0.7114910, 0.7717350, 0.0119784, 0.0897971, 0.2930210, 0.3238450, 0.8244310, 0.4989350, 0.9065360, 0.7243630, 0.6080610, 0.3995270, 0.7025980, 0.9413950, 0.4676490, 0.7364740, 0.9292950, 0.2833870, 0.7206830, 0.0787974, 0.7292470, 0.3833810, 0.9254370, 0.4232900, 0.3312770, 0.6945750, 0.1868070, 0.5928520, 0.9920520, 0.7017730, 0.1209040, 0.4473380, 0.7422080, 0.6688000, 0.9810240, 0.6444340, 0.2164730, 0.1661300, 0.0605885, 0.2900850, 0.9569210, 0.6231700, 0.8964550, 0.4904410, 0.1132310, 0.7994630, 0.0228514, 0.8074860, 0.3350700, 0.0078106, 0.6697860, 0.8061990, 0.9620900, 0.6584820, 0.9402010, 0.5316480, 0.4692150, 0.2955500, 0.8830100, 0.4025660, 0.9521750, 0.1921930, 0.7156490, 0.0509620, 0.5435290, 0.6958040, 0.5123500, 0.3825900, 0.9122690, 0.8171620, 0.1452080, 0.8154740, 0.0847717, 0.5643430, 0.4644440, 0.2725440, 0.4858110, 0.0429048, 0.8134510, 0.1922400, 0.4105230, 0.5632910, 0.4748170, 0.3086320, 0.4621590, 0.6638740, 0.3910020, 0.8894260, 0.6788130, 0.2051120, 0.6730940, 0.8837860, 0.0004909, 0.4109710, 0.3106920, 0.5159520, 0.7460340, 0.0091155, 0.3316360, 0.3155610, 0.4655370, 0.3144530, 0.8217770, 0.9635730, 0.9495410, 0.2787910, 0.1553760, 0.9618290, 0.8847550, 0.3721380, 0.2747430, 0.1392740, 0.9257780, 0.0532418, 0.7157340, 0.9172240, 0.6843300, 0.1728140, 0.5471560, 0.0285390, 0.3149070, 0.8884590, 0.6341110, 0.6789050, 0.3171770, 0.4468980, 0.4536390, 0.6995010, 0.3288150, 0.1677050, 0.3637050, 0.2355930, 0.3396380, 0.3991750, 0.9335000, 0.8455640, 0.9648870, 0.7714990, 0.5837530, 0.2914750, 0.5991130, 0.5860030, 0.6042740, 0.0678786, 0.7034880, 0.5017800, 0.2567860, 0.5917270, 0.3875160, 0.8740100, 0.5823080, 0.8106380, 0.3374130, 0.6663930, 0.7293340, 0.6518870, 0.8357480, 0.7972790, 0.2371150, 0.7593140, 0.9090090, 0.9780630, 0.5565970, 0.8128610, 0.0252937, 0.4484520, 0.5189970, 0.1129800, 0.6688300, 0.3643230, 0.3891070, 0.0650824, 0.7938640, 0.7312360, 0.7960090, 0.1902760, 0.7258130, 0.5245940, 0.9808760, 0.0645280, 0.6525940, 0.6528100, 0.3186540, 0.8609240, 0.5135930, 0.1139270, 0.8755680, 0.8149840, 0.5450900, 0.6120230, 0.9376900, 0.3170420, 0.2981590, 0.4241350, 0.8480880, 0.2283990, 0.5370940, 0.0093522, 0.0495578, 0.8347970, 0.8806240, 0.3195060, 0.5289380, 0.9454840, 0.7394620, 0.6555560, 0.4489600, 0.4819850, 0.8410490, 0.9721090, 0.9749600, 0.7500950, 0.8319440, 0.2599130, 0.2641030, 0.7377530, 0.7648360, 0.2238300, 0.9850640, 0.7085400, 0.1815490, 0.6203540, 0.5560750, 0.6541280, 0.5121810, 0.3872990, 0.6474720, 0.5936500, 0.1386580, 0.7985550, 0.5545780, 0.3958040, 0.7114390, 0.0268450, 0.0966318, 0.6370660, 0.9116560, 0.7222960, 0.5827630, 0.7240740, 0.0356666, 0.2560920, 0.7235860, 0.6229230, 0.0987210, 0.3529130, 0.4599630, 0.9366320, 0.1023150, 0.6442430, 0.5533250, 0.2779360, 0.7171610, 0.0069087, 0.6259890, 0.4710670, 0.8337760, 0.9197460, 0.2416770, 0.2671260, 0.2142710, 0.7875570, 0.2086330, 0.9999850, 0.6304560, 0.6027820, 0.2476110, 0.8080690, 0.7123560, 0.0063814, 0.6219940, 0.2666680, 0.6782140, 0.3568490, 0.5360430, 0.8681620, 0.4160270, 0.5564120, 0.6716780, 0.5991320, 0.5493000, 0.1838080, 0.9883280, 0.2243990, 0.3250140, 0.4686470, 0.7280790, 0.9565680, 0.9729910, 0.7638470, 0.7819340, 0.9977250, 0.5785990, 0.2603810, 0.1361900, 0.6748310, 0.7914580, 0.3620380, 0.8017590, 0.3533300, 0.1113830, 0.5578160, 0.2514450, 0.9703320, 0.3008020, 0.1695710, 0.6244220, 0.7367050, 0.6538350, 0.6229440, 0.4609500, 0.0458748, 0.1364850, 0.3836680, 0.2029540, 0.3383270, 0.1290850, 0.2096710, 0.9600260, 0.9683840, 0.5825560, 0.8090870, 0.4438490, 0.2991700, 0.0936808, 0.9771520, 0.0363587, 0.8494800, 0.5385000, 0.0298546, 0.3215480, 0.6589370, 0.6536010, 0.6138720, 0.6005790, 0.2702030, 0.6243300, 0.7878920, 0.4322420, 0.4292300, 0.9680100, 0.3775470, 0.0786398, 0.6516770, 0.3926360, 0.3841000, 0.8977920, 0.7522110, 0.1228160, 0.0022953, 0.6612420, 0.6404240, 0.6507160, 0.3557410, 0.7726500, 0.3489910, 0.2035280, 0.8672860, 0.2811420, 0.6150630, 0.9834950, 0.9078660, 0.2132660, 0.0484352, 0.4665030, 0.8185060, 0.3184980, 0.5529880, 0.0613801, 0.6795380, 0.9340690, 0.7692890, 0.9611750, 0.2030840, 0.8363350, 0.2945050, 0.7842040, 0.2851520, 0.1193780, 0.9128470, 0.0346805, 0.3525540, 0.2316420, 0.4011890, 0.4650280, 0.0865776, 0.7758880, 0.7430630, 0.9073090, 0.8585270, 0.7858130, 0.0447026, 0.9103100, 0.1666900, 0.7779020, 0.0135698, 0.4025940, 0.9675200, 0.3922060, 0.8357230, 0.5765260, 0.7672830, 0.4098370, 0.8333660, 0.7324780, 0.7818810, 0.2510220, 0.4681270, 0.5919410, 0.1856230, 0.9221090, 0.3411540, 0.5782570, 0.8058030, 0.6924370, 0.9798740, 0.0961788, 0.2020150, 0.0187089, 0.3036500, 0.1452400, 0.6908330, 0.9168720, 0.6539460, 0.5994230, 0.3231260, 0.8471000, 0.6657930, 0.3128600, 0.4755770, 0.8586220, 0.3377250, 0.6407820, 0.8242100, 0.0109879, 0.6323800, 0.0341605, 0.9882230, 0.6184880, 0.3310000, 0.7234350, 0.4325030, 0.2670900, 0.3881630, 0.7621760, 0.1780340, 0.5364270, 0.7759880, 0.2953840, 0.7000830, 0.6665840, 0.2929940, 0.5825120, 0.3788330, 0.7943280, 0.6663590, 0.9037930, 0.8053780, 0.6495870, 0.9443520, 0.8068080, 0.9374390, 0.9700780, 0.1335030, 0.5806630, 0.9737510, 0.3684750, 0.9747870, 0.5637450, 0.7599740, 0.2002640, 0.9933180, 0.4232000, 0.7824690, 0.1304800, 0.7678160, 0.5151630, 0.3876930, 0.6889290, 0.8225340, 0.7476470, 0.0253880, 0.7391240, 0.6938130, 0.2202260, 0.5404990, 0.8359890, 0.2912200, 0.6932400, 0.2344310, 0.0423549, 0.3640540, 0.8245590, 0.6384580, 0.3453230, 0.7002150, 0.7522460, 0.1580510, 0.3494370, 0.6230810, 0.6334450, 0.4055510, 0.4138450, 0.6761010, 0.5746230, 0.1597800, 0.6625530, 0.7055250, 0.3601730, 0.7777990, 0.0945425, 0.8528360, 0.0623906, 0.3733390, 0.0181806, 0.0900350, 0.5430030, 0.9535530, 0.4768050, 0.9385720, 0.5793960, 0.2177770, 0.6466360, 0.2385830, 0.6124740, 0.1378700, 0.6170460, 0.6187620, 0.3916250, 0.5590450, 0.4907770, 0.3549280, 0.2541050, 0.8260440, 0.2553220, 0.9594370, 0.9368440, 0.7658630, 0.0430100, 0.3356180, 0.7369050, 0.8216200, 0.9155720, 0.8995630, 0.4242420, 0.7547340, 0.3823430, 0.3504250, 0.1770410, 0.7962400, 0.0635463, 0.0081557, 0.1169980, 0.4546850, 0.1669870, 0.8784920, 0.8474790, 0.8791240, 0.4043130, 0.3932260, 0.1074270, 0.1946280, 0.0784943, 0.0243568, 0.2562060, 0.9510250, 0.8047630, 0.4923430, 0.7531020, 0.3965780, 0.9499460, 0.6503080, 0.7119420, 0.7861180, 0.5253750, 0.0496848, 0.6979340, 0.9649510, 0.1203280, 0.9826450, 0.7007020, 0.7201780, 0.5135590, 0.8317490, 0.3616720, 0.7505170, 0.0895694, 0.9106560, 0.7676280, 0.5551960, 0.4764760, 0.2676540, 0.0385173, 0.0407341, 0.6104580, 0.9861490, 0.1285120, 0.3513700, 0.9681440, 0.9317200, 0.9196610, 0.8307570, 0.1592440, 0.8678440, 0.1275210, 0.4027170, 0.2032900, 0.6260960, 0.2597440, 0.6135420, 0.0976725, 0.4993040, 0.4570500, 0.7663300, 0.4307250, 0.8635170, 0.4797700, 0.9090830, 0.7578530, 0.7851520, 0.7721210, 0.7233520, 0.4383730, 0.0651840, 0.7224350, 0.1688630, 0.8226180, 0.4175190, 0.1584690, 0.0435896, 0.7535050, 0.9365210, 0.0966345, 0.2711310, 0.7942350, 0.2504670, 0.7878460, 0.7332100, 0.9517010, 0.7224040, 0.5741370, 0.2665460, 0.8751080, 0.5013030, 0.5825900, 0.2271960, 0.5943400, 0.0316508, 0.4619630, 0.9864510, 0.5181610, 0.3797560, 0.7159930, 0.1677460, 0.3042100, 0.0220835, 0.7452070, 0.9591050, 0.6728300, 0.8024200, 0.8770700, 0.7300120, 0.3341970, 0.9278170, 0.1460310, 0.5898320, 0.1566060, 0.2215890, 0.0329922, 0.5396380, 0.7823650, 0.5524480, 0.5405200, 0.7242220, 0.2856190, 0.0056820, 0.8376220, 0.4172570, 0.7231610, 0.9057710, 0.6516550, 0.3143090, 0.8836300, 0.7463560, 0.3054240, 0.0774430, 0.3390590, 0.8778400, 0.4278040, 0.2951960, 0.7847920, 0.8547260, 0.6656660, 0.3087380, 0.9926950, 0.7833480, 0.2053050, 0.5043610, 0.8430290, 0.2443470, 0.7665600, 0.9709530, 0.5165540, 0.5897750, 0.9751420, 0.2774000, 0.6563290, 0.2604360, 0.6190380, 0.0912724, 0.1382830, 0.5270090, 0.4918650, 0.8638680, 0.6191290, 0.3426830, 0.1228050, 0.6938570, 0.6146970, 0.6679660, 0.7103110, 0.5653380, 0.5104620, 0.7145520, 0.5364350, 0.6699180, 0.3360010, 0.7718800, 0.0668492, 0.5731070, 0.7064920, 0.1220070, 0.5483620, 0.7825640, 0.9014250, 0.2072980, 0.1842920, 0.7006360, 0.6662320, 0.4618500, 0.0838058, 0.6726540, 0.6480640, 0.4279360, 0.6515050, 0.0100016, 0.1197710, 0.5707270, 0.1680100, 0.9809740, 0.4184610, 0.2763120, 0.3972900, 0.9552240, 0.6884780, 0.9711450, 0.6817630, 0.8360000, 0.3761510, 0.6317540, 0.7773180, 0.4952460, 0.8672210, 0.6982700, 0.8093750, 0.0612150, 0.2976580, 0.1909580, 0.7310600, 0.4555360, 0.6157010, 0.4223990, 0.0179701, 0.5192720, 0.5762930, 0.7454270, 0.1506500, 0.8256120, 0.9541790, 0.7986280, 0.5764040, 0.9627560, 0.4695920, 0.3707270, 0.7223370, 0.9990000, 0.0273482, 0.4021480, 0.1049750, 0.1857150, 0.5834740, 0.7794270, 0.5173930, 0.2450370, 0.8900850, 0.2008220, 0.9603760, 0.7406690, 0.9846990, 0.6642670, 0.3534440, 0.4286060, 0.2918950, 0.0034132, 0.3201140, 0.8712980, 0.7093740, 0.6984450, 0.0918986, 0.1741770, 0.9458920, 0.2720620, 0.7500820, 0.7621460, 0.2330300, 0.8666920, 0.5049790, 0.3562900, 0.7631770, 0.0749494, 0.6755260, 0.4509570, 0.3515390, 0.9399260, 0.9208810, 0.5356830, 0.5905670, 0.1931010, 0.0794843, 0.0264884, 0.6886080, 0.2469200, 0.7037440, 0.5908180, 0.5463110, 0.2490430, 0.4668820, 0.2645040, 0.9757230, 0.2363020, 0.0129618, 0.2680750, 0.6963430, 0.9530080, 0.8118140, 0.7405740, 0.5363450, 0.5889100, 0.0350188, 0.0539605, 0.8657040, 0.6226490, 0.6343820, 0.3438740, 0.1972660, 0.6592060, 0.3202850, 0.7464110, 0.7252530, 0.7901650, 0.5169400, 0.6057320, 0.1781070, 0.2226380, 0.8415510, 0.1341540, 0.3532300, 0.0445690, 0.7651240, 0.1124630, 0.3114470, 0.1770700, 0.4252710, 0.1282120, 0.5235500, 0.7107690, 0.9181580, 0.9655840, 0.5728210, 0.1677770, 0.9157200, 0.7763820, 0.6654540, 0.2381090, 0.8379170, 0.4007660, 0.3276580, 0.6526880, 0.1772620, 0.1836120, 0.5789990, 0.5513800, 0.0086409, 0.0059344, 0.5650960, 0.1686040, 0.0444728, 0.2203350, 0.2936010, 0.4379750, 0.0815387, 0.3875640, 0.6757950, 0.2464890, 0.9306980, 0.4755000, 0.0943825, 0.3629180, 0.3070490, 0.1845160, 0.2776860, 0.2683590, 0.5380870, 0.8239500, 0.6528460, 0.3367250, 0.6378520, 0.9281170, 0.7550990, 0.2171600, 0.9589480, 0.8821590, 0.1812970, 0.1039970, 0.6434080, 0.8452600, 0.6872650, 0.2299840, 0.5524580, 0.3595780, 0.4474590, 0.7775540, 0.5576080, 0.8446540, 0.4658620, 0.7817990, 0.5065020, 0.6282550, 0.9750010, 0.7155160, 0.5094850, 0.0134544, 0.9547380, 0.8664900, 0.0870459, 0.1962610, 0.8985950, 0.6893750, 0.6992920, 0.4354590, 0.5714150, 0.4448580, 0.8735020, 0.0501232, 0.0492682, 0.4518520, 0.2251710, 0.0703045, 0.2425590, 0.5553540, 0.7274430, 0.3289720, 0.1174910, 0.5384270, 0.1457230, 0.0518529, 0.1067330, 0.9649700, 0.6336400, 0.5407380, 0.2477960, 0.6949180, 0.3292640, 0.9465010, 0.8074960, 0.4773930, 0.2447020, 0.3745280, 0.0149108, 0.3947200, 0.8440610, 0.6580980, 0.4983170, 0.6294190, 0.4301880, 0.4766350, 0.1773510, 0.5951290, 0.8706510, 0.0415575, 0.7971230, 0.2770570, 0.5748970, 0.0126817, 0.1736770, 0.3195440, 0.1643600, 0.9692090, 0.2822370, 0.2570880, 0.7711970, 0.6102270, 0.1568450, 0.3963790, 0.7412440, 0.3831680, 0.2218230, 0.3073560, 0.0444407, 0.0335558, 0.7773800, 0.2444300, 0.0375941, 0.6234660, 0.4746180, 0.1802260, 0.8549260, 0.7781410, 0.9354720, 0.0394117, 0.4253140, 0.6244910, 0.0113432, 0.3984080, 0.6530700, 0.8472930, 0.7596740, 0.0896829, 0.9369430, 0.7380610, 0.7653090, 0.0963648, 0.6885130, 0.1974940, 0.3141560, 0.9870800, 0.8965770, 0.6767620, 0.3764350, 0.6673910, 0.2474220, 0.5390930, 0.1364230, 0.6236190, 0.0024082, 0.6977550, 0.2858700, 0.8603810, 0.5086290, 0.5626930, 0.5639980, 0.8966180, 0.1052880, 0.9275980, 0.4649430, 0.2175040, 0.5031210, 0.0068874, 0.2208880, 0.1668900, 0.1023200, 0.9050080, 0.1276970, 0.7688980, 0.9600920, 0.4892800, 0.2827210, 0.4446200, 0.6327600, 0.7488190, 0.0193288, 0.7328970, 0.1430370, 0.6839760, 0.6558340, 0.5708720, 0.1051340, 0.3381180, 0.8474480, 0.2693190, 0.8595110, 0.3836830, 0.7421180, 0.5815260, 0.6833340, 0.7375930, 0.1762440, 0.3290330, 0.7634410, 0.5607990, 0.3324150, 0.5279050, 0.3850710, 0.4301150, 0.8124000, 0.9911360, 0.6035760, 0.1856210, 0.1638350, 0.9970130, 0.4125290, 0.7650510, 0.7742160, 0.4228200, 0.7762360, 0.0043048, 0.4681560, 0.5772460, 0.7725860, 0.1948970, 0.0427962, 0.8289050, 0.0889241, 0.3405560, 0.3822820, 0.0470675, 0.0724488, 0.1278800, 0.7361160, 0.9816510, 0.8783470, 0.7220060, 0.3551090, 0.8164350, 0.9978180, 0.8404960, 0.4081490, 0.7703870, 0.4315360, 0.7692100, 0.6545580, 0.9536040, 0.6320800, 0.7142060, 0.3565320, 0.3559030, 0.4631340, 0.4746390, 0.9884300, 0.2920340, 0.2063970, 0.1119370, 0.3031480, 0.0495715, 0.1871950, 0.3082640, 0.8626140, 0.4568540, 0.7531260, 0.6847490, 0.6160270, 0.4936120, 0.9389500, 0.6879530, 0.5596080, 0.7911590, 0.5139580, 0.9674970, 0.3947800, 0.4991370, 0.8523360, 0.8464800, 0.6474510, 0.6351240, 0.7704790, 0.4332760, 0.9302390, 0.7752350, 0.6860520, 0.0721703, 0.1039230, 0.7858640, 0.5887420, 0.4709910, 0.3530540, 0.4260530, 0.1158660, 0.5504900, 0.1986780, 0.3433900, 0.2700010, 0.9151670, 0.1606500, 0.4011430, 0.4763370, 0.3125030, 0.1292500, 0.7530150, 0.8208750, 0.2598140, 0.4689550, 0.4310740, 0.7855690, 0.1384650, 0.6926870, 0.2236260, 0.8043500, 0.6812940, 0.5541100, 0.7024750, 0.9520530, 0.7545800, 0.2319930, 0.5054190, 0.8941920, 0.4772430, 0.1249770, 0.7011860, 0.1475100, 0.3164740, 0.5319350, 0.9548490, 0.8034350, 0.7159960, 0.8069010, 0.7665480, 0.6665960, 0.5511290, 0.3354490, 0.6906760, 0.1308100, 0.6676750, 0.0911185, 0.8097650, 0.0010914, 0.7168160, 0.7814880, 0.2531780, 0.3458810, 0.7337600, 0.5685250, 0.3764640, 0.6995190, 0.8535620, 0.8054270, 0.2624120, 0.4265180, 0.3278870, 0.0923758, 0.0878845, 0.3745980, 0.9477080, 0.0973729, 0.8588640, 0.2769770, 0.8759400, 0.4261670, 0.1516060, 0.4016950, 0.0569647, 0.2820340, 0.4472430, 0.0252490, 0.1040980, 0.2254310, 0.4764620, 0.6984700, 0.9571160, 0.2305970, 0.3931590, 0.1130070, 0.1872240, 0.4622620, 0.5619620, 0.7887350, 0.6344100, 0.8203910, 0.2022090, 0.7392210, 0.8257760, 0.8812100, 0.7308220, 0.7251490, 0.2503480, 0.9252280, 0.8120080, 0.4216130, 0.3126680, 0.7898050, 0.1095550, 0.7856660, 0.5756690, 0.2943090, 0.9977590, 0.7502660, 0.4771040, 0.0611894, 0.7956290, 0.6237990, 0.0964943, 0.6992220, 0.0874087, 0.1472820, 0.0475997, 0.2912380, 0.3821950, 0.1396160, 0.3097380, 0.0651353, 0.5712570, 0.9858860, 0.2951240, 0.0333507, 0.6649520, 0.8612090, 0.1842190, 0.3770160, 0.0818375, 0.7852160, 0.0088950, 0.2603340, 0.7983110, 0.6251010, 0.9970280, 0.1603900, 0.7318280, 0.7619560, 0.7841730, 0.8085100, 0.6765670, 0.1559590, 0.8713950, 0.7364920, 0.0281426, 0.9654640, 0.8164060, 0.1284310, 0.8984070, 0.5726220, 0.5946100, 0.8369550, 0.5897960, 0.6526580, 0.7779090, 0.5360280, 0.5217690, 0.9920650, 0.8056090, 0.6735180, 0.1301100, 0.3212450, 0.0459818, 0.8617790, 0.5539260, 0.4366310, 0.7973430, 0.7169120, 0.1773760, 0.2208730, 0.9051140, 0.6667640, 0.9774600, 0.8141700, 0.4351820, 0.6478940, 0.1692750, 0.7520330, 0.5375520, 0.7445940, 0.1887650, 0.2410040, 0.9262390, 0.5764870, 0.0603974, 0.2677450, 0.4516830, 0.6973320, 0.5428710, 0.1626230, 0.9369350, 0.8825160, 0.6520220, 0.9449710, 0.9795960, 0.2616590, 0.1232150, 0.2046530, 0.7712620, 0.9245190, 0.2526570, 0.9578050, 0.0609674, 0.8485200, 0.2112200, 0.9889020, 0.4603020, 0.4399450, 0.0630004, 0.9099480, 0.7223610, 0.3228370, 0.4084820, 0.1049020, 0.0407128, 0.9019170, 0.2828360, 0.5233480, 0.2740490, 0.3415380, 0.7594860, 0.7628130, 0.0723421, 0.3165420, 0.0468863, 0.3582200, 0.8941540, 0.7938160, 0.0945285, 0.9634730, 0.6415240, 0.7623290, 0.7685580, 0.0711655, 0.0663946, 0.7865980, 0.2497690, 0.6764170, 0.4335670, 0.9268590, 0.8938080, 0.2687750, 0.2211010, 0.7394210, 0.6686800, 0.7700900, 0.7216010, 0.6312810, 0.3851290, 0.7484730, 0.3617550, 0.0844655, 0.5118940, 0.5191290, 0.9348060, 0.3164320, 0.5142220, 0.8965020, 0.8879330, 0.5373510, 0.0193262, 0.0045669, 0.8178890, 0.9623230, 0.4053250, 0.3570500, 0.4113530, 0.7396370, 0.3099780, 0.7748530, 0.0121860, 0.8558350, 0.9488930, 0.5341490, 0.4596180, 0.5681150, 0.5048890, 0.5685400, 0.5645450, 0.4115280, 0.7663360, 0.3928310, 0.8280610, 0.2251540, 0.1310120, 0.6826810, 0.2502480, 0.0069636, 0.8647690, 0.4028470, 0.8727550, 0.3326970, 0.5226970, 0.0687790, 0.7391630, 0.8094370, 0.9275760, 0.9223230, 0.7189840, 0.9135360, 0.7791080, 0.6281690, 0.7609960, 0.2844840, 0.4374700, 0.3194420, 0.3640480, 0.6782890, 0.6221670, 0.0718088, 0.5155360, 0.9936200, 0.5380980, 0.6678080, 0.6335250, 0.3895570, 0.0780268, 0.2950020, 0.0253779, 0.7866260, 0.9974990, 0.1083550, 0.7793400, 0.6918410, 0.5308120, 0.9250680, 0.4372120, 0.1746830, 0.2107390, 0.9580150, 0.1077090, 0.7690700, 0.9409440, 0.2617820, 0.6909020, 0.5468840, 0.1678840, 0.3596560, 0.5880960, 0.9414020, 0.2743980, 0.2004320, 0.8707950, 0.7525440, 0.0837463, 0.6830420, 0.4061220, 0.1279520, 0.3651580, 0.9611160, 0.0478651, 0.6589560, 0.0258810, 0.4396360, 0.1029980, 0.7675420, 0.4166460, 0.2820690, 0.8086060, 0.3877760, 0.8788420, 0.2970440, 0.1012890, 0.2035720, 0.1404780, 0.7885790, 0.1982100, 0.3214810, 0.7621580, 0.6010150, 0.7642950, 0.7092050, 0.1785810, 0.6166120, 0.0514721, 0.7280450, 0.6084110, 0.7478640, 0.3900680, 0.5793850, 0.5901040, 0.9569530, 0.3071500, 0.7662830, 0.0685652, 0.5132400, 0.9145130, 0.8490610, 0.3024670, 0.7351470, 0.6090060, 0.6982600, 0.9503760, 0.5519360, 0.5423930, 0.7804410, 0.1913170, 0.9259370, 0.3857550, 0.0165344, 0.2379340, 0.1813710, 0.1043760, 0.6721550, 0.4756910, 0.4030690, 0.9300050, 0.1532780, 0.2989340, 0.6553250, 0.9136410, 0.3741250, 0.1133450, 0.6171610, 0.0209665, 0.0784943, 0.1168410, 0.0356596, 0.7405910, 0.9451200, 0.6597330, 0.0175239, 0.8763220, 0.3257870, 0.7105260, 0.7391460, 0.0923020, 0.0868425, 0.7775350, 0.6980800, 0.8416590, 0.8788010, 0.4829710, 0.4372180, 0.6452400, 0.3743250, 0.6024750, 0.6903570, 0.7446300, 0.4440690, 0.0478554, 0.0923863, 0.1772160, 0.7713310, 0.2814190, 0.9969390, 0.8825890, 0.6430500, 0.0730902, 0.2970940, 0.4383160, 0.9199670, 0.8809470, 0.5680600, 0.0259789, 0.7655180, 0.4934100, 0.7223920, 0.1453460, 0.2343760, 0.0785597, 0.4923920, 0.3928540, 0.2221090, 0.6750910, 0.3389080, 0.4138160, 0.8514940, 0.9462430, 0.0719682, 0.1439420, 0.7551590, 0.4466590, 0.8551780, 0.0207658, 0.5066330, 0.8672430, 0.4539870, 0.8590780, 0.9588840, 0.0746826, 0.2623220, 0.3003070, 0.3599200, 0.0145316, 0.4655430, 0.3883140, 0.6050470, 0.4075390, 0.5454620, 0.2595910, 0.1476760, 0.6046500, 0.7621070, 0.2934070, 0.7020250, 0.1342610, 0.1776630, 0.3463120, 0.5996590, 0.6093580, 0.6413450, 0.2615290, 0.1453490, 0.5059500, 0.4156580, 0.7678470, 0.4803070, 0.1634970, 0.2265040, 0.8759050, 0.0873939, 0.6663450, 0.6209800, 0.5578770, 0.1977560, 0.7615140, 0.1786520, 0.0149915, 0.3428780, 0.0566734, 0.7038380, 0.9774340, 0.2240760, 0.1544050, 0.4177380, 0.5478810, 0.5194950, 0.7423760, 0.6509550, 0.2098790, 0.4357940, 0.8141130, 0.3239710, 0.9471490, 0.3241850, 0.1893210, 0.5841120, 0.7138880, 0.5506460, 0.3271790, 0.1574240, 0.4197220, 0.5084220, 0.4101050, 0.0257217, 0.0129424, 0.0174187, 0.8622440, 0.3414990, 0.9025160, 0.3336980, 0.9701990, 0.5423520, 0.0708323, 0.0385804, 0.6426330, 0.4291600, 0.3285560, 0.5001660, 0.9464210, 0.5104530, 0.9735040, 0.3726420, 0.5843330, 0.9765840, 0.2659090, 0.0046825, 0.8658210, 0.2727080, 0.5871870, 0.8348930, 0.9117290, 0.2509300, 0.1119530, 0.4046500, 0.0533098, 0.4369620, 0.0776575, 0.3785200, 0.9500030, 0.1645810, 0.5654370, 0.2655560, 0.9682200, 0.7141250, 0.7051070, 0.1198060, 0.9594930, 0.4427160, 0.3300100, 0.9048680, 0.6163820, 0.6741360, 0.1462050, 0.2061420, 0.2446880, 0.3900730, 0.5980900, 0.1472150, 0.9907220, 0.1117660, 0.7574110, 0.8656740, 0.3022400, 0.7581890, 0.9659730, 0.4105600, 0.4845310, 0.0280272, 0.3181180, 0.2854710, 0.6748080, 0.3360900, 0.0225539, 0.8911060, 0.2541100, 0.6270100, 0.7377010, 0.0071696, 0.8359210, 0.7372730, 0.1792090, 0.3216730, 0.8721970, 0.1516150, 0.8819450, 0.2163450, 0.8433530, 0.8680000, 0.0915683, 0.0258308, 0.6309370, 0.1800680, 0.2280030, 0.9081640, 0.1310990, 0.8766490, 0.0029961, 0.2465370, 0.8380300, 0.5050910, 0.2413550, 0.2013100, 0.1973770, 0.7653590, 0.5961430, 0.7433650, 0.2133840, 0.4350530, 0.2205770, 0.7762280, 0.2138340, 0.8661220, 0.3890340, 0.1095670, 0.0464561, 0.0832056, 0.3997330, 0.0262677, 0.4029120, 0.8395370, 0.4669670, 0.4398140, 0.8262910, 0.1013930, 0.0951412, 0.2059460, 0.7638540, 0.5586080, 0.4618410, 0.7370140, 0.7884620, 0.9654640, 0.6252450, 0.3757040, 0.8109070, 0.1237050, 0.8556310, 0.6344930, 0.7971080, 0.3548940, 0.8722950, 0.4507720, 0.3652980, 0.0512534, 0.8754080, 0.5194120, 0.1762830, 0.7764710, 0.5454500, 0.1611470, 0.2827400, 0.9496750, 0.0152315, 0.9018850, 0.7657170, 0.5916640, 0.1275490, 0.4290510, 0.7298050, 0.3080710, 0.4270940, 0.6701920, 0.2295540, 0.1441090, 0.1330210, 0.6216070, 0.8465130, 0.5029560, 0.3359140, 0.1323340, 0.6592770, 0.3355220, 0.7135750, 0.9413530, 0.0011651, 0.5061080, 0.6118750, 0.5149220, 0.0172299, 0.7299520, 0.4506250, 0.4392480, 0.7239140, 0.2123710, 0.0552749, 0.1894100, 0.0994915, 0.1257220, 0.2107280, 0.8141840, 0.5488930, 0.4292660, 0.0916592, 0.5846920, 0.8841030, 0.3634590, 0.8866060, 0.9161480, 0.9878600, 0.0438769, 0.8450390, 0.5130790, 0.3832450, 0.1706040, 0.5913760, 0.7773790, 0.1514520, 0.6758090, 0.3018510, 0.8232460, 0.3103450, 0.0529507, 0.1995370, 0.2551330, 0.3589260, 0.2483630, 0.2839030, 0.1493840, 0.0457304, 0.1301510, 0.1592020, 0.4789420, 0.0136515, 0.2712260, 0.6050190, 0.7686170, 0.4895670, 0.0866235, 0.1113490, 0.5233270, 0.9996760, 0.9401910, 0.4462570, 0.4856430, 0.3535740, 0.5580960, 0.7425350, 0.7235610, 0.6404330, 0.7055770, 0.9348210, 0.8191290, 0.4305680, 0.0915904, 0.2608620, 0.6461380, 0.8226030, 0.3465350, 0.7042570, 0.5767130, 0.8055990, 0.2478780, 0.7023260, 0.3508710, 0.8013230, 0.1179540, 0.4020030, 0.4992880, 0.7853330, 0.7451510, 0.4696930, 0.3652010, 0.1253540, 0.1434870, 0.8592910, 0.0702645, 0.0031832, 0.0092401, 0.7294880, 0.3808060, 0.0670584, 0.6458100, 0.7278110, 0.6735030, 0.8124350, 0.9895220, 0.9223200, 0.2625160, 0.0829659, 0.0608477, 0.7011200, 0.7665310, 0.6554390, 0.8131830, 0.2799770, 0.5577760, 0.5779560, 0.0002941, 0.8624740, 0.4095410, 0.5419870, 0.9652020, 0.9547510, 0.9105580, 0.1570910, 0.6574070, 0.7227620, 0.8958820, 0.4605000, 0.9217780, 0.2471380, 0.0443455, 0.4271960, 0.7032110, 0.8217430, 0.3511870, 0.2873590, 0.6609190, 0.8895120, 0.9819960, 0.1363570, 0.9239850, 0.0641371, 0.2835010, 0.4286840, 0.2842750, 0.6104190, 0.0371339, 0.4820110, 0.2223960, 0.4792200, 0.2223910, 0.7407010, 0.0931516, 0.1414630, 0.5615480, 0.7445230, 0.1165210, 0.5007720, 0.9821480, 0.0353092, 0.9822340, 0.5982690, 0.5793110, 0.1682290, 0.8933760, 0.4496080, 0.5038680, 0.7111840, 0.9090110, 0.5756770, 0.8575070, 0.3185830, 0.8481950, 0.5885000, 0.4637900, 0.6428070, 0.0770022, 0.7106920, 0.6698550, 0.9009440, 0.5507390, 0.8923480, 0.1957240, 0.7600680, 0.4575700, 0.3686740, 0.1067320, 0.2578920, 0.4835720, 0.6635970, 0.7559700, 0.8002770, 0.8406960, 0.3886140, 0.3317160, 0.0373206, 0.5136170, 0.4517790, 0.5282280, 0.1321790, 0.3226850, 0.7965250, 0.6188380, 0.4488470, 0.8999440, 0.5745400, 0.5516340, 0.1387910, 0.5323340, 0.6336960, 0.0458351, 0.7682370, 0.6755560, 0.5729540, 0.8886120, 0.2531270, 0.5359110, 0.2994880, 0.1750150, 0.3331190, 0.4183800, 0.1638600, 0.5635680, 0.9141380, 0.3631030, 0.0262723, 0.2620550, 0.4382060, 0.8534020, 0.9511270, 0.2887200, 0.9933290, 0.2916990, 0.4552610, 0.1876130, 0.1836180, 0.7604600, 0.1969480, 0.9525840, 0.1437670, 0.5907120, 0.7248490, 0.5654090, 0.2997110, 0.2770750, 0.3710660, 0.9115440, 0.6613320, 0.3211230, 0.1463330, 0.6802970, 0.7996280, 0.2138150, 0.2878030, 0.6542010, 0.9770760, 0.9957250, 0.1230360, 0.0390928, 0.6840200, 0.5635730, 0.6070990, 0.2559600, 0.7766060, 0.0170484, 0.0929866, 0.1931890, 0.6425620, 0.9558150, 0.3814000, 0.1964340, 0.6097390, 0.6192180, 0.5251030, 0.0715810, 0.5421060, 0.1910190, 0.4364860, 0.6268040, 0.7637290, 0.6651430, 0.5972270, 0.4367380, 0.4280200, 0.9902360, 0.8941410, 0.8492340, 0.0850443, 0.5860530, 0.1319110, 0.0455448, 0.3274160, 0.6575320, 0.6382460, 0.6241710, 0.0768733, 0.1867280, 0.3091940, 0.1994010, 0.9570790, 0.8310600, 0.7954600, 0.6057230, 0.3766210, 0.9168270, 0.1092400, 0.3692830, 0.3483540, 0.3669010, 0.1184520, 0.3034890, 0.0012791, 0.2608630, 0.4923940, 0.8680300, 0.2784520, 0.1245520, 0.6719730, 0.1802380, 0.8085390, 0.7848490, 0.4676010, 0.4209640, 0.3422220, 0.8485730, 0.3992010, 0.7968580, 0.7495290, 0.7148030, 0.4488270, 0.7529000, 0.7018720, 0.9189580, 0.2665000, 0.6539900, 0.4402900, 0.6931850, 0.2807440, 0.1113070, 0.5903140, 0.2923770, 0.4997840, 0.9507870, 0.7922690, 0.1605550, 0.7016930, 0.9192710, 0.1722300, 0.7350430, 0.9667770, 0.6750530, 0.6902620, 0.8243980, 0.2231760, 0.1964580, 0.6448440, 0.3766920, 0.2979010, 0.9969990, 0.2411830, 0.1461740, 0.8466140, 0.8711600, 0.5767870, 0.1176920, 0.3256100, 0.5606520, 0.5404030, 0.4767010, 0.6917630, 0.8839050, 0.4797870, 0.3273020, 0.4907160, 0.7885520, 0.0644317, 0.3341610, 0.4869960, 0.5692780, 0.8609170, 0.3233210, 0.7188390, 0.6394630, 0.4065270, 0.2902470, 0.2607390, 0.1527280, 0.9035660, 0.4056590, 0.1350190, 0.1786280, 0.0695994, 0.3599140, 0.8688660, 0.7084580, 0.6430070, 0.2380460, 0.7388280, 0.9675340, 0.5190410, 0.2072280, 0.4059390, 0.4201900, 0.2852580, 0.2269050, 0.4873070, 0.8721030, 0.2442900, 0.0018687, 0.1272650, 0.1168260, 0.4302490, 0.1341680, 0.7968840, 0.9425920, 0.3618100, 0.3574830, 0.9748300, 0.9287740, 0.2202030, 0.1595630, 0.4187440, 0.2199730, 0.4022430, 0.7254200, 0.0133862, 0.4553320, 0.9211430, 0.3677670, 0.6842960, 0.3460760, 0.7271880, 0.6530610, 0.8457060, 0.8958200, 0.3379870, 0.3546130, 0.5119520, 0.1477830, 0.2853390, 0.0165682, 0.7179650, 0.8446680, 0.9998220, 0.9319990, 0.9475600, 0.9651930, 0.2056540, 0.2916510, 0.4198170, 0.3933410, 0.6103600, 0.1765250, 0.3172300, 0.7301380, 0.9415000, 0.9466870, 0.9982460, 0.2074430, 0.8673770, 0.6537060, 0.2521350, 0.4532190, 0.1701890, 0.9484420, 0.3427300, 0.1908050, 0.2544490, 0.3381430, 0.1676560, 0.5876710, 0.8213210, 0.9850870, 0.5614910, 0.7822640, 0.8194700, 0.1277530, 0.3304980, 0.4699970, 0.8623620, 0.2994320, 0.1173460, 0.8709460, 0.9093270, 0.3533130, 0.7273040, 0.7052160, 0.4661910, 0.9589010, 0.8934450, 0.8371680, 0.8480890, 0.8863180, 0.3245010, 0.2386070, 0.9473030, 0.5004300, 0.9700990, 0.7842490, 0.9493430, 0.5388960, 0.1873010, 0.9057350, 0.5785130, 0.1980810, 0.3064830, 0.0313068, 0.8679730, 0.6303110, 0.1746320, 0.2251780, 0.2142350, 0.7214970, 0.1656840, 0.8044540, 0.2690470, 0.0576627, 0.8277390, 0.3094160, 0.2493910, 0.2830920, 0.8721940, 0.2533480, 0.9680800, 0.3245930, 0.6720680, 0.9813140, 0.1065300, 0.1396620, 0.6265390, 0.7018760, 0.5745100, 0.8556170, 0.7126500, 0.0795662, 0.3664850, 0.1114670, 0.6797190, 0.2302240, 0.1717060, 0.8639860, 0.0001290, 0.1381140, 0.7617410, 0.6740780, 0.5975560, 0.8206830, 0.7245780, 0.9903880, 0.6024690, 0.6267230, 0.5722730, 0.0176668, 0.0912659, 0.1048180, 0.1246580, 0.9674200, 0.8287320, 0.4055210, 0.6290040, 0.3985850, 0.9521790, 0.1038620, 0.9230050, 0.7226460, 0.8583690, 0.4027690, 0.7559350, 0.7419370, 0.9682780, 0.3802990, 0.1565250, 0.3831730, 0.3221670, 0.9705970, 0.4041600, 0.6308200, 0.1278890, 0.7669760, 0.7231030, 0.5005480, 0.8274040, 0.3967540, 0.1273580, 0.6391740, 0.5115590, 0.2390260, 0.0773237, 0.5718770, 0.0417843, 0.6018310, 0.4800090, 0.0834750, 0.0511570, 0.8449930, 0.2949830, 0.6131190, 0.8586430, 0.6818160, 0.3665460, 0.7695900, 0.0068255, 0.9467400, 0.4777820, 0.3157900, 0.6063660, 0.2089570, 0.6825690, 0.4196930, 0.3691370, 0.5261380, 0.1221880, 0.3818510, 0.2715950, 0.0502835, 0.5787870, 0.5531360, 0.5641530, 0.8149370, 0.4743310, 0.8073240, 0.9362880, 0.8514270, 0.3200110, 0.9348860, 0.4886780, 0.9225200, 0.9518480, 0.3315700, 0.6974720, 0.7020880, 0.2956450, 0.7249110, 0.5230120, 0.9434010, 0.3922210, 0.2428310, 0.3054780, 0.1667330, 0.0132527, 0.2106360, 0.5641590, 0.4783690, 0.7643060, 0.2162800, 0.6916660, 0.9723200, 0.5622700, 0.4371630, 0.8337700, 0.3823460, 0.5614670, 0.0855501, 0.5032710, 0.3014790, 0.2612470, 0.6218230, 0.8311780, 0.9577290, 0.1288050, 0.2181710, 0.1331840, 0.0423000, 0.5338720, 0.6420350, 0.2122880, 0.8777150, 0.8277780, 0.4033820, 0.7009840, 0.2520720, 0.3643210, 0.1421930, 0.6776560, 0.3743710, 0.1999880, 0.4679990, 0.1192090, 0.9847850, 0.6009100, 0.6533140, 0.8595030, 0.7020820, 0.0005596, 0.4049150, 0.6647960, 0.3249660, 0.1784550, 0.6384680, 0.0991271, 0.6593460, 0.9688290, 0.1396820, 0.9230800, 0.2886110, 0.8721840, 0.4792390, 0.9838460, 0.1020230, 0.8576370, 0.8071740, 0.0976768, 0.5284340, 0.4054190, 0.7235720, 0.9547470, 0.6690990, 0.4348070, 0.8114950, 0.1965430, 0.7286010, 0.8812620, 0.7949660, 0.6659530, 0.0850262, 0.9189380, 0.9525500, 0.5774210, 0.9547300, 0.0729483, 0.7285060, 0.4013470, 0.9738890, 0.4468910, 0.7882430, 0.3971950, 0.4053680, 0.2679620, 0.0007739, 0.6031570, 0.5302070, 0.6396310, 0.2331250, 0.1459950, 0.8053220, 0.6287560, 0.3971460, 0.2925540, 0.3566160, 0.3475990, 0.0258548, 0.7650200, 0.2816160, 0.5909210, 0.4554700, 0.9839010, 0.3437200, 0.0822885, 0.4059500, 0.1315080, 0.7500430, 0.1062350, 0.1205720, 0.0239533, 0.9499170, 0.1012160, 0.0050358, 0.4658790, 0.4418090, 0.8994590, 0.3547680, 0.6142060, 0.6764890, 0.3675380, 0.5214740, 0.5642910, 0.4442210, 0.7994220, 0.1397500, 0.8284060, 0.2026190, 0.6655360, 0.9786060, 0.7676450, 0.9409070, 0.2664950, 0.6817710, 0.7640920, 0.4408890, 0.3350920, 0.2856680, 0.6589110, 0.9167360, 0.1442920, 0.1697180, 0.2143000, 0.2150880, 0.1892620, 0.0219648, 0.9866160, 0.4867280, 0.1611680, 0.2495050, 0.4462110, 0.8573510, 0.5606500, 0.3307360, 0.3636190, 0.1621730, 0.9032090, 0.4094850, 0.2369730, 0.5226120, 0.5204420, 0.4406470, 0.5274730, 0.2546360, 0.9427170, 0.9839020, 0.4279480, 0.9584410, 0.6671470, 0.3180260, 0.0084008, 0.2488500, 0.6186170, 0.7822630, 0.7131310, 0.9859930, 0.3435060, 0.2132350, 0.4624290, 0.9577050, 0.2214680, 0.4484430, 0.6419870, 0.2832540, 0.6395330, 0.6400830, 0.1236860, 0.0550310, 0.1410670, 0.0707865, 0.8018600, 0.3524930, 0.4057450, 0.6299450, 0.8080200, 0.7364140, 0.7221320, 0.5335980, 0.3284500, 0.7346290, 0.2833950, 0.3667530, 0.6396080, 0.5837020, 0.2915190, 0.5894730, 0.4546220, 0.7772300, 0.6712160, 0.3062140, 0.8501810, 0.9443080, 0.6451050, 0.2886940, 0.6250880, 0.0026797, 0.3559000, 0.4302860, 0.4967410, 0.8028160, 0.5441120, 0.8692590, 0.5996270, 0.7768950, 0.7899830, 0.1117140, 0.0474378, 0.5071840, 0.8508200, 0.4734870, 0.8965690, 0.5026650, 0.0744139, 0.8246260, 0.7117330, 0.7586210, 0.2285370, 0.0276296, 0.6342030, 0.6799020, 0.8293590, 0.8488960, 0.4434070, 0.2811540, 0.6563070, 0.7176330, 0.5547630, 0.8218910, 0.1689120, 0.9364460, 0.0254215, 0.8674760, 0.0609941, 0.2645770, 0.9066640, 0.5775310, 0.6719890, 0.8779100, 0.1892170, 0.3977930, 0.8308460, 0.7689650, 0.0512993, 0.3555090, 0.6132600, 0.2991190, 0.5563710, 0.7488830, 0.6977620, 0.5981930, 0.2014560, 0.6573180, 0.8159660, 0.8789530, 0.6857870, 0.8259550, 0.3836320, 0.1022620, 0.1823970, 0.2521290, 0.4693440, 0.3635580, 0.5747370, 0.6247940, 0.1436100, 0.0573465, 0.3125890, 0.5500810, 0.5733280, 0.3966010, 0.5242500, 0.5495050, 0.8183870, 0.5539960, 0.7073840, 0.5926380, 0.5617530, 0.6574390, 0.1015850, 0.5384860, 0.1445060, 0.5870780, 0.2939730, 0.8714550, 0.3475720, 0.9050160, 0.2328190, 0.7941750, 0.8986020, 0.8115840, 0.0961899, 0.4750300, 0.7609390, 0.3610130, 0.4724500, 0.4182470, 0.8626870, 0.9681770, 0.5420570, 0.2304710, 0.2918370, 0.2121030, 0.0880626, 0.6535620, 0.8356420, 0.0965102, 0.8540730, 0.4259790, 0.0560160, 0.0084900, 0.2554090, 0.2614460, 0.5049640, 0.8256070, 0.2959120, 0.1573390, 0.5460140, 0.3867390, 0.9303740, 0.7608870, 0.7728100, 0.4571830, 0.4702560, 0.3681430, 0.2243810, 0.2307190, 0.1104250, 0.0836710, 0.8499340, 0.3059980, 0.5399300, 0.6279510, 0.4277030, 0.1499160, 0.6138620, 0.1201330, 0.2480650, 0.0833317, 0.5022360, 0.0876848, 0.0203285, 0.0594994, 0.6044050, 0.6498630, 0.3338470, 0.9742630, 0.6157180, 0.3360600, 0.8861210, 0.7210360, 0.1876410, 0.2155950, 0.2663720, 0.9120710, 0.6774410, 0.3656770, 0.5639500, 0.2613830, 0.6302150, 0.7861810, 0.6469350, 0.9559310, 0.5344610, 0.9553740, 0.8900800, 0.8414450, 0.2569390, 0.1499240, 0.0443634, 0.1562060, 0.2279290, 0.5598240, 0.1373450, 0.1091300, 0.0820987, 0.3072970, 0.5114090, 0.2849060, 0.2917410, 0.1317710, 0.3461720, 0.5958060, 0.6718260, 0.4483460, 0.8118540, 0.5230230, 0.6871880, 0.8473250, 0.0019612, 0.1977720, 0.9146870, 0.4804080, 0.9518620, 0.4032180, 0.2142530, 0.2994380, 0.5372510, 0.8682230, 0.4849760, 0.3894700, 0.5589550, 0.3402890, 0.3929080, 0.0800373, 0.9815020, 0.3694010, 0.7891410, 0.2692750, 0.8968790, 0.2855440, 0.4308070, 0.4481670, 0.8329470, 0.8360970, 0.5801280, 0.6177140, 0.7821190, 0.8272320, 0.6223300, 0.7613110, 0.7047840, 0.0675711, 0.3884710, 0.1647600, 0.0705471, 0.9500470, 0.8123890, 0.4698630, 0.7746840, 0.5079670, 0.1218390, 0.8183870, 0.0410639, 0.5962130, 0.1447850, 0.2039340, 0.3614490, 0.0603859, 0.4565000, 0.3336370, 0.3997030, 0.5019520, 0.5112190, 0.8398540, 0.0163766, 0.4788320, 0.2446000, 0.3335860, 0.4040950, 0.9819780, 0.7417710, 0.3132670, 0.4105230, 0.5862100, 0.5306080, 0.6359890, 0.9139010, 0.9578820, 0.1364750, 0.7507810, 0.0971772, 0.1598730, 0.4285160, 0.7123820, 0.9645260, 0.0601257, 0.8968020, 0.2792430, 0.5477930, 0.4153830, 0.7692190, 0.2734100, 0.1022450, 0.9857940, 0.4797910, 0.2081600, 0.1631230, 0.2802000, 0.4902910, 0.7783200, 0.2210280, 0.2537370, 0.4938840, 0.3494830, 0.1081080, 0.7408420, 0.6065550, 0.1764460, 0.7360290, 0.3313550, 0.8091510, 0.6397890, 0.2934900, 0.5917720, 0.1644430, 0.3301010, 0.2725450, 0.1417350, 0.0428891, 0.6710680, 0.9949180, 0.2612030, 0.6156770, 0.8702780, 0.1319980, 0.5282880, 0.3975950, 0.2357770, 0.2055020, 0.7693810, 0.2330350, 0.8083630, 0.5600380, 0.5294560, 0.0702819, 0.0874801, 0.0855406, 0.2778640, 0.3977970, 0.0761266, 0.7308080, 0.6802340, 0.3429650, 0.1897030, 0.5383870, 0.3047650, 0.0349436, 0.7779730, 0.7727340, 0.4636920, 0.5327770, 0.3996770, 0.4657820, 0.8281060, 0.0360405, 0.7857590, 0.9327050, 0.8654120, 0.2803900, 0.6662230, 0.3323770, 0.2733620, 0.3961650, 0.6761550, 0.5872550, 0.9746770, 0.4011590, 0.7823650, 0.1328940, 0.0017993, 0.0980254, 0.3473810, 0.1496390, 0.8161820, 0.4645070, 0.1910060, 0.3066330, 0.9208290, 0.7360620, 0.4384970, 0.5709180, 0.4618800, 0.1920920, 0.3021170, 0.4011780, 0.0460099, 0.7686840, 0.5225510, 0.1158060, 0.9866030, 0.5673300, 0.8590460, 0.4749980, 0.8179880, 0.3433620, 0.0886746, 0.9212200, 0.0816793, 0.5042290, 0.8243290, 0.0129333, 0.6558210, 0.1135380, 0.5436680, 0.7675370, 0.5786570, 0.0970849, 0.0914784, 0.8392460, 0.5445640, 0.1214740, 0.8769040, 0.0959044, 0.9324830, 0.3388370, 0.9709230, 0.5117980, 0.8810830, 0.2103990, 0.0956102, 0.8305970, 0.7942270, 0.0840216, 0.7672350, 0.8149750, 0.4783640, 0.2406060, 0.2498330, 0.2775760, 0.9458990, 0.4343200, 0.7820760, 0.9522200, 0.9500210, 0.2597320, 0.3015720, 0.1396730, 0.2912260, 0.1016880, 0.5991610, 0.4721570, 0.2143830, 0.4746200, 0.6991570, 0.5461910, 0.5093950, 0.3480720, 0.4905330, 0.1306100, 0.7968670, 0.8677100, 0.8521760, 0.4107360, 0.7982130, 0.7174220, 0.7672900, 0.9772710, 0.6027350, 0.1408490, 0.6937350, 0.9011750, 0.3601170, 0.6733080, 0.6877230, 0.2035930, 0.8265470, 0.9684160, 0.7187410, 0.4613680, 0.3058870, 0.4635830, 0.9826290, 0.6359460, 0.3482400, 0.8009380, 0.5037560, 0.8181410, 0.9451060, 0.1799380, 0.3132620, 0.0942642, 0.0882643, 0.1079410, 0.7821690, 0.2842140, 0.0575928, 0.3004970, 0.9930920, 0.3091630, 0.6821140, 0.3254680, 0.6620430, 0.8598350, 0.6051430, 0.9939090, 0.0486293, 0.4518140, 0.6817250, 0.7701910, 0.8144840, 0.3481350, 0.2337220, 0.4526470, 0.7703850, 0.4155850, 0.3565220, 0.4620780, 0.3973520, 0.0061075, 0.3479110, 0.8148620, 0.8032280, 0.3965930, 0.5485910, 0.1252560, 0.4995200, 0.3625450, 0.9789950, 0.2659280, 0.5378290, 0.3398540, 0.9502100, 0.5370130, 0.1125110, 0.5724170, 0.7613620, 0.9599190, 0.2215330, 0.8330590, 0.5226970, 0.6692390, 0.4480040, 0.4986270, 0.2856670, 0.8385550, 0.6522670, 0.5319600, 0.1131320, 0.6317170, 0.0255143, 0.5676720, 0.3005730, 0.3280110, 0.2498060, 0.5565840, 0.1328870, 0.7569580, 0.8287750, 0.0632252, 0.9968670, 0.7404920, 0.1936450, 0.2996780, 0.1638610, 0.8013690, 0.0076874, 0.3882780, 0.1253470, 0.0600926, 0.3474680, 0.3601980, 0.8581750, 0.4651690, 0.2123560, 0.9176480, 0.0251175, 0.5613700, 0.9012700, 0.0422091, 0.9064570, 0.2647890, 0.9214960, 0.4226440, 0.1153640, 0.9862440, 0.2280650, 0.0862243, 0.3527750, 0.4601270, 0.8132220, 0.0280067, 0.6449600, 0.2965800, 0.2965640, 0.6771770, 0.5000680, 0.9825050, 0.1244910, 0.9799450, 0.5314270, 0.3128220, 0.3238520, 0.1330740, 0.4864170, 0.4745110, 0.5574350, 0.5291260, 0.1879120, 0.4945290, 0.2652980, 0.9276720, 0.2094500, 0.1435330, 0.8876060, 0.2892010, 0.3627350, 0.0225607, 0.5343460, 0.7899290, 0.9465130, 0.0447000, 0.7406690, 0.4986760, 0.7197040, 0.4004310, 0.0162218, 0.2379240, 0.9342810, 0.1863440, 0.5957560, 0.8160340, 0.1020330, 0.9445410, 0.6752530, 0.9387000, 0.0284920, 0.1072290, 0.9635100, 0.1924620, 0.9751720, 0.9292160, 0.6653770, 0.0700025, 0.8369320, 0.7796600, 0.0476228, 0.3886690, 0.0504397, 0.8029670, 0.6056680, 0.6574350, 0.9604670, 0.1173790, 0.0497091, 0.0918100, 0.7689140, 0.3547710, 0.9330440, 0.5593710, 0.3398760, 0.6504000, 0.6251280, 0.3371830, 0.5868900, 0.6977930, 0.6063370, 0.8247690, 0.3670850, 0.0153332, 0.2360320, 0.0973758, 0.5894850, 0.4480980, 0.0148679, 0.4287720, 0.2056950, 0.8314030, 0.4816650, 0.3664470, 0.0533304, 0.6563510, 0.9225130, 0.6240390, 0.2951950, 0.0679228, 0.1501290, 0.5923930, 0.8031130, 0.7329940, 0.7135250, 0.7039760, 0.8782710, 0.6188160, 0.7897490, 0.3722440, 0.4439940, 0.7503160, 0.1812870, 0.6790020, 0.3744300, 0.3121040, 0.1155030, 0.1268760, 0.3393310, 0.9178600, 0.9514670, 0.4658360, 0.6443180, 0.6277640, 0.1503880, 0.0208179, 0.6063190, 0.0381839, 0.1879980, 0.4859850, 0.9207910, 0.1035740, 0.1203730, 0.9564030, 0.8837750, 0.1223640, 0.7708280, 0.4987160, 0.3569410, 0.2987490, 0.5012630, 0.1702670, 0.3103180, 0.3708550, 0.2696690, 0.3562720, 0.2682230, 0.3557650, 0.5786020, 0.9485850, 0.5036550, 0.9294470, 0.4959340, 0.8793730, 0.3906160, 0.8383060, 0.6484730, 0.0466035, 0.9876450, 0.2972020, 0.2926860, 0.1874760, 0.7323850, 0.1570090, 0.0118404, 0.4170510, 0.9195160, 0.5380540, 0.1532130, 0.3706150, 0.4441170, 0.7702260, 0.9370070, 0.6289950, 0.2770950, 0.9267470, 0.1519030, 0.9164490, 0.4089000, 0.7244510, 0.6102800, 0.4079650, 0.6726440, 0.5230490, 0.5616390, 0.1480780, 0.1172700, 0.6733610, 0.8468800, 0.7811890, 0.6480000, 0.1534570, 0.3893470, 0.8259310, 0.2282180, 0.2445270, 0.1101670, 0.6901570, 0.1751240, 0.6806910, 0.0253786, 0.5509380, 0.3660090, 0.1591900, 0.1612420, 0.7736780, 0.5954390, 0.8221410, 0.5888830, 0.7693730, 0.2572730, 0.4718840, 0.0551648, 0.6995290, 0.7253010, 0.8096890, 0.9439640, 0.4908170, 0.2876750, 0.6784840, 0.7122910, 0.7446120, 0.7354240, 0.7781700, 0.0302992, 0.6857280, 0.0426081, 0.0082657, 0.6265690, 0.1397490, 0.1904440, 0.3984140, 0.5058150, 0.1100890, 0.7094600, 0.0826661, 0.6023670, 0.7626170, 0.0984021, 0.6628460, 0.7523860, 0.2693520, 0.9850760, 0.5758090, 0.7306980, 0.3143910, 0.3361110, 0.0499767, 0.2867330, 0.3018220, 0.1317790, 0.6861780, 0.3951560, 0.0037069, 0.1615980, 0.6197000, 0.3772080, 0.3667770, 0.2491750, 0.6611090, 0.3920470, 0.6211160, 0.6187980, 0.1391870, 0.5498120, 0.3834160, 0.7267770, 0.6355550, 0.2175970, 0.4686270, 0.1084600, 0.5759540, 0.3285840, 0.5885920, 0.8025820, 0.8814370, 0.6036050, 0.6108000, 0.2068490, 0.0696173, 0.7047130, 0.5998490, 0.4088820, 0.2391000, 0.4276860, 0.0656017, 0.6347140, 0.4871570, 0.4769660, 0.9471110, 0.2987940, 0.9183190, 0.0077897, 0.2901390, 0.1621810, 0.6472530, 0.9207050, 0.8038150, 0.0791085, 0.0830087, 0.7793180, 0.6407350, 0.1474220, 0.7131370, 0.6743470, 0.5367850, 0.0082303, 0.2450870, 0.2305850, 0.0109471, 0.1968250, 0.4834710, 0.9328600, 0.4943040, 0.3001380, 0.9551380, 0.6654750, 0.7424260, 0.5216130, 0.6303110, 0.8661050, 0.7503180, 0.2910490, 0.5890560, 0.4015950, 0.2566230, 0.9637210, 0.8781100, 0.2292600, 0.1893760, 0.1225010, 0.7762930, 0.9669650, 0.1960980, 0.7794550, 0.0278145, 0.0407415, 0.8958140, 0.1568590, 0.9471880, 0.8723790, 0.2402770, 0.5580650, 0.2964970, 0.9755750, 0.3959650, 0.8579740, 0.4504520, 0.7801960, 0.1744590, 0.2253850, 0.8939780, 0.8831380, 0.5382660, 0.6592420, 0.9932700, 0.7441050, 0.6121640, 0.1390790, 0.6307220, 0.3852540, 0.1384530, 0.9997140, 0.6492930, 0.8855640, 0.4877290, 0.9125830, 0.6586500, 0.5444390, 0.4095000, 0.3350550, 0.7647030, 0.1645830, 0.1093370, 0.4928860, 0.4998690, 0.7602550, 0.8710610, 0.0542912, 0.5817210, 0.5029060, 0.4332070, 0.8662580, 0.5985070, 0.5339190, 0.3234320, 0.4919120, 0.8808520, 0.0238407, 0.9987790, 0.7612670, 0.7762150, 0.7368510, 0.3710980, 0.1732650, 0.1675210, 0.4074470, 0.7376080, 0.6382160, 0.9883340, 0.5213350, 0.2173770, 0.1854180, 0.7449600, 0.6458840, 0.7814160, 0.6082940, 0.2960940, 0.2565430, 0.1701950, 0.9441500, 0.8704380, 0.0413776, 0.4663530, 0.4814380, 0.3245210, 0.4071870, 0.7238910, 0.3025310, 0.5773060, 0.8970340, 0.6032290, 0.8019760, 0.6331210, 0.6790910, 0.7316060, 0.5249810, 0.2343630, 0.6957210, 0.1999800, 0.7288720, 0.7795850, 0.2491560, 0.0539375, 0.5189060, 0.7243860, 0.5725550, 0.1905330, 0.7624550, 0.6284980, 0.6761320, 0.8827390, 0.8895560, 0.8994920, 0.6533910, 0.0420752, 0.5559590, 0.7495140, 0.4158780, 0.3770090, 0.8968400, 0.5025900, 0.2418730, 0.3459380, 0.7998610, 0.7632110, 0.8007430, 0.0030635, 0.0101395, 0.4930200, 0.5179170, 0.4599700, 0.6348220, 0.4372340, 0.8826020, 0.1375400, 0.9383770, 0.0017237, 0.3832010, 0.9461780, 0.0604190, 0.6892610, 0.8432520, 0.5198000, 0.2168390, 0.1250040, 0.6401070, 0.6140970, 0.8213300, 0.7870640, 0.2115800, 0.7063930, 0.9752020, 0.1227730, 0.0876060, 0.2141120, 0.1354870, 0.2024670, 0.3695880, 0.2666480, 0.1386320, 0.2599790, 0.9964630, 0.7048400, 0.1670200, 0.6357640, 0.9973200, 0.0968092, 0.8688110, 0.7262780, 0.7980620, 0.6653790, 0.5460360, 0.4146530, 0.8923790, 0.3590460, 0.1648410, 0.3894550, 0.8408680, 0.7345860, 0.3129540, 0.6196670, 0.6302120, 0.6918640, 0.1522600, 0.6842670, 0.2554400, 0.2855310, 0.7513870, 0.4988360, 0.1786620, 0.2733180, 0.4898150, 0.5011110, 0.1577590, 0.7380220, 0.4707420, 0.4705190, 0.3810870, 0.3835810, 0.9858420, 0.1636620, 0.6236180, 0.8964400, 0.3011510, 0.2637920, 0.1082870, 0.7437180, 0.4899330, 0.2648030, 0.1211690, 0.9266950, 0.3968800, 0.3198890, 0.8415370, 0.6061290, 0.8362660, 0.1204590, 0.3217660, 0.2927570, 0.7236980, 0.8824520, 0.8631910, 0.6957310, 0.9919430, 0.8018760, 0.0647500, 0.3730150, 0.4947460, 0.8884090, 0.4847940, 0.9424140, 0.8144660, 0.6491170, 0.9723620, 0.0550595, 0.3391330, 0.0373841, 0.1884230, 0.4865080, 0.2771230, 0.4173210, 0.9033010, 0.1362290, 0.8455110, 0.5932800, 0.8142260, 0.0467882, 0.0024829, 0.5865610, 0.7204870, 0.6174070, 0.2873020, 0.3235500, 0.7923760, 0.6716160, 0.8233970, 0.5017480, 0.3889970, 0.0155549, 0.0983678, 0.0255883, 0.3859270, 0.3521500, 0.6906610, 0.7409280, 0.9973510, 0.6743850, 0.5520020, 0.3769820, 0.5894490, 0.7914430, 0.2957740, 0.3734790, 0.9938200, 0.0284342, 0.9153160, 0.8546140, 0.6574000, 0.9072990, 0.8472480, 0.9983620, 0.1007720, 0.0324397, 0.2040840, 0.8839330, 0.9829900, 0.9057130, 0.8678370, 0.1416300, 0.7224180, 0.9091480, 0.6633530, 0.2210870, 0.6859600, 0.8544320, 0.1101630, 0.8826820, 0.8408830, 0.8066620, 0.2366200, 0.0586061, 0.2396210, 0.2498300, 0.0945670, 0.9309130, 0.0131086, 0.3998460, 0.0264227, 0.2889190, 0.3812630, 0.8595860, 0.8562780, 0.1935000, 0.5255820, 0.3488370, 0.8061540, 0.4033900, 0.4842330, 0.1839340, 0.1018630, 0.4707080, 0.4662660, 0.2909130, 0.4338740, 0.8112380, 0.8058840, 0.9422270, 0.6297100, 0.1033790, 0.6997970, 0.7101160, 0.0558575, 0.0871777, 0.3599200, 0.1466920, 0.4919070, 0.3321330, 0.3138160, 0.0268018, 0.4627930, 0.3821020, 0.2759340, 0.4272220, 0.9195850, 0.3801280, 0.1501650, 0.7313650, 0.0134822, 0.7138760, 0.4593620, 0.8986920, 0.7420370, 0.1450520, 0.0410450, 0.3176300, 0.0446820, 0.3639390, 0.5987090, 0.6015850, 0.0563388, 0.4481410, 0.5911490, 0.2868260, 0.8565220, 0.0007120, 0.1478030, 0.7715820, 0.6508800, 0.2725070, 0.3027970, 0.8533170, 0.1833250, 0.6347190, 0.8379430, 0.4222280, 0.5506090, 0.1866210, 0.1410440, 0.0562423, 0.5048990, 0.5817590, 0.2116510, 0.2496570, 0.3701700, 0.3644420, 0.8089070, 0.2188300, 0.7153080, 0.7170640, 0.3246970, 0.6263090, 0.5578900, 0.0351741, 0.0209612, 0.6986790, 0.3388950, 0.5088530, 0.9367020, 0.7793640, 0.8862290, 0.0587639, 0.1464790, 0.1536930, 0.1211680, 0.7522820, 0.2484230, 0.8792620, 0.4302480, 0.7276300, 0.6280450, 0.0539065, 0.5360970, 0.9384220, 0.6430280, 0.0259859, 0.8768050, 0.6784270, 0.9303030, 0.4543840, 0.3833150, 0.6581090, 0.4684950, 0.1018970, 0.6053600, 0.3656860, 0.8297570, 0.0283219, 0.7727060, 0.3442660, 0.0806821, 0.2749690, 0.2954090, 0.3690000, 0.1748020, 0.5861910, 0.5325600, 0.8067490, 0.2560880, 0.6812820, 0.6137460, 0.9100600, 0.4145200, 0.8000290, 0.4064900, 0.9076480, 0.1147730, 0.4058960, 0.1525050, 0.6482850, 0.8846130, 0.1969610, 0.0505325, 0.9500130, 0.0607249, 0.5845630, 0.8752860, 0.9669670, 0.0998430, 0.8881510, 0.4983070, 0.0334989, 0.7905040, 0.9138290, 0.5211990, 0.4066300, 0.8838810, 0.0858788, 0.7945010, 0.6708330, 0.2343390, 0.5720410, 0.2118720, 0.2412420, 0.3491640, 0.2561140, 0.9936360, 0.1447500, 0.6987310, 0.2098880, 0.5224660, 0.0802735, 0.1932780, 0.8566730, 0.6319790, 0.3321740, 0.7954950, 0.5589260, 0.5834740, 0.6435640, 0.6858320, 0.7088790, 0.9464660, 0.9527540, 0.8134340, 0.9903650, 0.9981210, 0.6555360, 0.3689700, 0.9199030, 0.7575050, 0.1119100, 0.3947380, 0.8155910, 0.9285370, 0.3798750, 0.6087240, 0.0492550, 0.3108640, 0.9334790, 0.9655590, 0.2272510, 0.7965230, 0.6460080, 0.6204780, 0.2489830, 0.7341630, 0.3940680, 0.7482310, 0.4233180, 0.6640530, 0.7186390, 0.6001000, 0.8102060, 0.1111010, 0.5781420, 0.7586650, 0.9160740, 0.6526340, 0.9058880, 0.9014560, 0.3518630, 0.1927210, 0.3333140, 0.3091160, 0.6527850, 0.5315540, 0.5908510, 0.3570710, 0.5490960, 0.1059330, 0.7831660, 0.5168510, 0.8674390, 0.3923530, 0.0169184, 0.7923330, 0.3881210, 0.7497220, 0.7454970, 0.7263480, 0.4268400, 0.3647150, 0.2375530, 0.4307700, 0.9510850, 0.1129180, 0.6275320, 0.9447370, 0.5998860, 0.8074550, 0.1338310, 0.5337300, 0.7422330, 0.4503900, 0.3648980, 0.3082920, 0.2907020, 0.2206810, 0.1131310, 0.4866600, 0.7445360, 0.7004850, 0.7287680, 0.0245126, 0.1406730, 0.2314660, 0.4473880, 0.9088960, 0.4642250, 0.9214180, 0.8515140, 0.6987630, 0.6018500, 0.7386590, 0.6356690, 0.7188160, 0.8381000, 0.1688720, 0.7086460, 0.8565360, 0.6871640, 0.1354780, 0.3919200, 0.2664070, 0.3230500, 0.5391090, 0.6344450, 0.3645520, 0.9693690, 0.7248950, 0.9756050, 0.2874620, 0.3915920, 0.6595900, 0.3611000, 0.6881290, 0.4123920, 0.7807400, 0.4412640, 0.3505320, 0.7660160, 0.1863450, 0.1505670, 0.2040490, 0.3092740, 0.0461331, 0.0947103, 0.8275810, 0.8798250, 0.7893630, 0.9566940, 0.7667840, 0.1052410, 0.2986460, 0.4611000, 0.5770380, 0.8288600, 0.2272650, 0.3276020, 0.0796657, 0.8877560, 0.1019260, 0.2284830, 0.4033830, 0.6284000, 0.3556370, 0.3107630, 0.2824850, 0.8494750, 0.4310940, 0.8381730, 0.3339620, 0.3859450, 0.3603180, 0.0402893, 0.2467810, 0.5434580, 0.6704780, 0.9923830, 0.6899600, 0.9500730, 0.1531590, 0.3654170, 0.6021250, 0.0909522, 0.5762480, 0.6056010, 0.6871650, 0.9200180, 0.6477240, 0.8310770, 0.5079340, 0.9963730, 0.7247490, 0.7005140, 0.2955740, 0.6503570, 0.9068400, 0.9424110, 0.9897860, 0.6227540, 0.4585510, 0.1207700, 0.8585380, 0.6251090, 0.2713850, 0.7128310, 0.4678390, 0.4348960, 0.5448140, 0.3526450, 0.1154430, 0.8378710, 0.7072210, 0.2455120, 0.7399790, 0.5195180, 0.8957540, 0.5848530, 0.9933790, 0.3176420, 0.5754530, 0.3665580, 0.3031230, 0.1073560, 0.9894950, 0.2461590, 0.4235090, 0.2543680, 0.3924580, 0.1433370, 0.1401990, 0.5998510, 0.1359460, 0.9469980, 0.2795160, 0.8712260, 0.6408330, 0.1368370, 0.9240770, 0.8537870, 0.1218870, 0.7789590, 0.3306210, 0.3260980, 0.6903050, 0.6163520, 0.6426680, 0.6455580, 0.8896320, 0.6290700, 0.2323400, 0.0786784, 0.9686900, 0.7762500, 0.8466490, 0.7545900, 0.4110550, 0.0073691, 0.9346070, 0.9066450, 0.0239874, 0.6946570, 0.9742290, 0.0131753, 0.1546910, 0.0891958, 0.1231460, 0.8037910, 0.5485770, 0.3299780, 0.5633020, 0.7334950, 0.7819890, 0.8740120, 0.0975398, 0.7879230, 0.2000720, 0.9021510, 0.8294260, 0.1309380, 0.0963207, 0.8663340, 0.2072120, 0.7468900, 0.0892845, 0.7975900, 0.4209790, 0.8510410, 0.6902640, 0.1339740, 0.0138155, 0.7855840, 0.2024030, 0.5282130, 0.7564800, 0.3802920, 0.7743960, 0.0835906, 0.4464210, 0.8672790, 0.6792640, 0.4461360, 0.0588798, 0.1891070, 0.2929200, 0.4094360, 0.2977020, 0.7689140, 0.3426840, 0.5247920, 0.8280830, 0.1555140, 0.5590720, 0.9465190, 0.8357740, 0.3618790, 0.6632140, 0.8766460, 0.0203786, 0.8223060, 0.6116040, 0.6274070, 0.4477680, 0.7135110, 0.4995740, 0.0725222, 0.3950960, 0.7008780, 0.5682960, 0.5961690, 0.2522210, 0.9671790, 0.8892580, 0.4202720, 0.7110560, 0.8214100, 0.3086810, 0.9906890, 0.0030521, 0.3415230, 0.3442150, 0.4919600, 0.3568920, 0.9762040, 0.3370840, 0.8615730, 0.1248880, 0.7441730, 0.6087860, 0.4114860, 0.0283545, 0.6804440, 0.7838560, 0.5821960, 0.2539770, 0.2443970, 0.3939950, 0.4635070, 0.3602430, 0.0276459, 0.5802500, 0.4714680, 0.9016160, 0.2602580, 0.4472150, 0.5994950, 0.6892700, 0.1864470, 0.0920067, 0.4583410, 0.8082310, 0.9164860, 0.6892970, 0.1846950, 0.9890430, 0.1597550, 0.1490470, 0.3185200, 0.3694070, 0.2093430, 0.5273420, 0.1829290, 0.0220162, 0.1497760, 0.4399650, 0.3706940, 0.6723170, 0.1078350, 0.8470280, 0.5361400, 0.9595930, 0.5426830, 0.1687790, 0.9570260, 0.1405360, 0.9816910, 0.4046200, 0.2102520, 0.6550210, 0.4013920, 0.8394080, 0.4290990, 0.9761170, 0.0174025, 0.1568600, 0.2677660, 0.3611680, 0.1793100, 0.1138040, 0.9295890, 0.4823750, 0.9716340, 0.6777510, 0.8252760, 0.1395690, 0.0659684, 0.1892250, 0.1667030, 0.8546460, 0.8132990, 0.4779200, 0.8658910, 0.8963830, 0.7743760, 0.4886470, 0.3518740, 0.3787520, 0.1933230, 0.2227220, 0.0623922, 0.9063680, 0.0406616, 0.1716850, 0.5084030, 0.0704672, 0.9342890, 0.3194950, 0.4015450, 0.3084860, 0.8499580, 0.4550380, 0.7819910, 0.8470630, 0.9846530, 0.4978420, 0.6548620, 0.9428640, 0.9307670, 0.8422630, 0.6667980, 0.1510560, 0.9123730, 0.0745303, 0.3538460, 0.3441860, 0.5141510, 0.5927870, 0.6255520, 0.1939610, 0.7700660, 0.5806560, 0.8909450, 0.3806840, 0.6191150, 0.9520130, 0.8626860, 0.1349940, 0.3902490, 0.5912050, 0.1405520, 0.3976320, 0.2103880, 0.6073920, 0.0858505, 0.0414652, 0.4968270, 0.6039280, 0.9994540, 0.7412660, 0.1830000, 0.6152630, 0.8977470, 0.2112230, 0.4802590, 0.1939030, 0.7935990, 0.6773330, 0.1473230, 0.0436061, 0.7290120, 0.3787100, 0.2249100, 0.2124720, 0.4918050, 0.8627460, 0.6909480, 0.4115210, 0.2507250, 0.2351320, 0.1171670, 0.0063103, 0.8502750, 0.6656300, 0.2273930, 0.7820410, 0.4213920, 0.7937250, 0.3358990, 0.7482300, 0.6874030, 0.6275550, 0.9641520, 0.2086590, 0.6631410, 0.1873200, 0.0927388, 0.1058460, 0.3386750, 0.3238320, 0.8781280, 0.6715510, 0.6004140, 0.7407430, 0.2520590, 0.0838138, 0.2540690, 0.8912930, 0.6996810, 0.9125860, 0.1661610, 0.6269840, 0.0690349, 0.8440420, 0.5954250, 0.2854620, 0.2723570, 0.8308800, 0.5952660, 0.3467850, 0.0057564, 0.7157700, 0.6894270, 0.4697210, 0.5973720, 0.6256150, 0.8521120, 0.9351440, 0.0373541, 0.7920510, 0.7630950, 0.9474100, 0.8542990, 0.1603100, 0.4097390, 0.7030590, 0.3196540, 0.3771570, 0.4532500, 0.6165670, 0.9245190, 0.0248657, 0.5517660, 0.0994327, 0.8813170, 0.9957440, 0.9661430, 0.0613026, 0.6871310, 0.6115230, 0.6302710, 0.5618310, 0.2373920, 0.0948762, 0.2763510, 0.3773150, 0.6514290, 0.2535480, 0.5694080, 0.8108260, 0.2998410, 0.0941780, 0.6369510, 0.3562710, 0.9771440, 0.2501350, 0.8934150, 0.2218200, 0.0965918, 0.1329990, 0.0412172, 0.2311700, 0.7863410, 0.8212450, 0.8572490, 0.2855170, 0.2538670, 0.6184560, 0.9370770, 0.6350780, 0.2574060, 0.6848500, 0.1498630, 0.1664260, 0.5835640, 0.2590900, 0.3928190, 0.9248720, 0.0748873, 0.8802840, 0.0466396, 0.3679970, 0.2407880, 0.0319334, 0.7072740, 0.7812050, 0.8474740, 0.8646240, 0.4055760, 0.0266453, 0.4376760, 0.4178160, 0.6770090, 0.4320400, 0.0269236, 0.9095520, 0.3440810, 0.5108790, 0.1167910, 0.0582152, 0.2435480, 0.2135390, 0.5498640, 0.6067360, 0.8111940, 0.1660360, 0.9611420, 0.6176650, 0.3114670, 0.6873880, 0.8181560, 0.6140060, 0.5975080, 0.1563550, 0.6984530, 0.5965160, 0.7752930, 0.8015810, 0.9355500, 0.1028330, 0.8143080, 0.9153580, 0.9449910, 0.3310640, 0.7643620, 0.9786050, 0.0354411, 0.4272660, 0.6555990, 0.5813310, 0.6150630, 0.6202160, 0.4568420, 0.7110150, 0.1219990, 0.5779300, 0.2735340, 0.3701850, 0.7017150, 0.1851780, 0.8648990, 0.9156250, 0.6503320, 0.7568350, 0.2960740, 0.6337780, 0.2218300, 0.9896850, 0.5207130, 0.2660910, 0.9925580, 0.8773630, 0.5746930, 0.4445990, 0.5077260, 0.6353910, 0.5923270, 0.0199489, 0.5369900, 0.7580870, 0.6390090, 0.6964630, 0.0963926, 0.3287880, 0.1800410, 0.2400200, 0.2825940, 0.2369160, 0.8800370, 0.2609500, 0.4136930, 0.6102260, 0.9259710, 0.1464540, 0.3079720, 0.4097220, 0.4812360, 0.5149000, 0.3438780, 0.2224960, 0.7701270, 0.6397660, 0.8350850, 0.0336279, 0.7813200, 0.7826800, 0.2066410, 0.9398250, 0.1806710, 0.1549940, 0.1759450, 0.8629280, 0.1725180, 0.5518000, 0.8619370, 0.5091160, 0.6309030, 0.7243470, 0.5685870, 0.3355310, 0.7841530, 0.3382360, 0.3963540, 0.9289450, 0.9618190, 0.9951920, 0.7085110, 0.1623120, 0.0063451, 0.1242470, 0.8200880, 0.3034740, 0.6533570, 0.3006900, 0.6216270, 0.3999680, 0.0646744, 0.2991100, 0.0911747, 0.9408580, 0.6627920, 0.2296500, 0.5578730, 0.8105820, 0.2899300, 0.1684210, 0.4917260, 0.1027670, 0.6946530, 0.8962410, 0.0094068, 0.0447834, 0.1145370, 0.3132710, 0.0239673, 0.2114270, 0.2095430, 0.1482140, 0.2605220, 0.3044290, 0.5005300, 0.0722659, 0.0418213, 0.5871220, 0.0966995, 0.5918560, 0.9360860, 0.9696860, 0.5104390, 0.8622330, 0.9013960, 0.2275700, 0.9588060, 0.4251770, 0.1059510, 0.9408710, 0.0882869, 0.2933980, 0.1424260, 0.3468320, 0.8400450, 0.5592450, 0.1900100, 0.8153660, 0.5905390, 0.2182870, 0.9985860, 0.6081420, 0.6956120, 0.5935370, 0.1000070, 0.2067160, 0.1868700, 0.0571705, 0.8911060, 0.6333100, 0.6374300, 0.2088130, 0.2998000, 0.1590380, 0.7587570, 0.2240970, 0.8349290, 0.2335350, 0.1638050, 0.9204570, 0.4407720, 0.4886760, 0.9597540, 0.4586790, 0.7619430, 0.7005010, 0.4451210, 0.9514190, 0.8566540, 0.4843870, 0.6386360, 0.7970120, 0.7483460, 0.3180270, 0.0208344, 0.5033710, 0.8482360, 0.7191790, 0.7050640, 0.3562650, 0.4385050, 0.0102155, 0.0657357, 0.7171810, 0.5950540, 0.9625360, 0.3331530, 0.9207490, 0.7539180, 0.9136620, 0.6079410, 0.9892130, 0.6159460, 0.0252931, 0.8903980, 0.4649350, 0.7422440, 0.5582940, 0.1680840, 0.2427340, 0.1335140, 0.0425172, 0.0040355, 0.4138000, 0.8915480, 0.2275040, 0.6364580, 0.0250353, 0.2987050, 0.9721190, 0.6215070, 0.9731980, 0.3169250, 0.4301640, 0.6369370, 0.4455860, 0.3247050, 0.5777780, 0.9263240, 0.4082880, 0.0188897, 0.6743960, 0.6891530, 0.8195230, 0.3250620, 0.1218980, 0.1388050, 0.3332870, 0.5421430, 0.0157072, 0.7816860, 0.5021210, 0.0752774, 0.1542930, 0.0773440, 0.3779300, 0.5652450, 0.2313660, 0.7805280, 0.0406983, 0.3526080, 0.6259210, 0.6862620, 0.8525800, 0.7080590, 0.6053410, 0.5429840, 0.6379170, 0.4517960, 0.3203740, 0.6436580, 0.4987020, 0.0958287, 0.6758000, 0.5491110, 0.1055130, 0.5450930, 0.8411260, 0.7644380, 0.4145130, 0.2774140, 0.2605300, 0.5981380, 0.3164560, 0.0820851, 0.7511730, 0.9361680, 0.5960560, 0.2800140, 0.7253330, 0.3361330, 0.3464370, 0.9203510, 0.7740150, 0.7093800, 0.7042900, 0.4767890, 0.3615760, 0.4676640, 0.9058520, 0.2366580, 0.9903110, 0.1169940, 0.6372200, 0.3525470, 0.2739270, 0.4768170, 0.1863610, 0.0243964, 0.9542310, 0.8101560, 0.7120160, 0.0403057, 0.5504480, 0.4901500, 0.2794450, 0.7305570, 0.1669830, 0.3396080, 0.6611960, 0.1390770, 0.7621020, 0.5088990, 0.3935470, 0.8396740, 0.6968370, 0.4087610, 0.6150570, 0.7182380, 0.3882350, 0.0600654, 0.7375680, 0.8750870, 0.0263838, 0.8912190, 0.7778700, 0.8795880, 0.7684900, 0.3054980, 0.6403390, 0.4666000, 0.4495640, 0.6340420, 0.9748360, 0.7356210, 0.1065130, 0.1889770, 0.5627760, 0.7945520, 0.4560840, 0.8676420, 0.2450200, 0.1532100, 0.3400500, 0.8666070, 0.3580980, 0.9354260, 0.5720310, 0.5479540, 0.4465200, 0.0719223, 0.4427410, 0.0558807, 0.8871810, 0.6399010, 0.0037945, 0.2672200, 0.1949800, 0.1645210, 0.1527430, 0.6281470, 0.2232550, 0.3286960, 0.9777740, 0.1617290, 0.9222390, 0.2496360, 0.7941450, 0.4681000, 0.4436850, 0.9954490, 0.5275960, 0.2032520, 0.4186430, 0.7032250, 0.2024300, 0.1713900, 0.2809390, 0.2527280, 0.0851798, 0.7938800, 0.1580700, 0.7344060, 0.4911950, 0.7238390, 0.3366510, 0.1683910, 0.0915661, 0.2584910, 0.3402430, 0.9889300, 0.6331820, 0.1298190, 0.1617020, 0.3175460, 0.9788770, 0.1972070, 0.2165700, 0.2723490, 0.3353210, 0.8818310, 0.5626950, 0.2991310, 0.8929840, 0.4653620, 0.2288530, 0.2996760, 0.4791970, 0.1964750, 0.2559190, 0.8891600, 0.0652560, 0.2915620, 0.7560310, 0.8005680, 0.7622130, 0.1391650, 0.9730070, 0.5119410, 0.5484770, 0.2383390, 0.9175710, 0.2807010, 0.3462100, 0.9676420, 0.1812350, 0.9682070, 0.4566410, 0.6380830, 0.8725350, 0.9806890, 0.7664520, 0.3001220, 0.4098940, 0.1099500, 0.2458550, 0.4965100, 0.2609060, 0.1046770, 0.2970370, 0.8282500, 0.5353760, 0.9086930, 0.3882740, 0.4230860, 0.2355230, 0.9871260, 0.8024460, 0.2405950, 0.9608170, 0.3994630, 0.9837470, 0.4961530, 0.1378450, 0.7220410, 0.4847740, 0.5166330, 0.5506260, 0.0707650, 0.6236600, 0.7664830, 0.2714970, 0.9052200, 0.7474420, 0.4675210, 0.5675520, 0.5792030, 0.3894780, 0.9707870, 0.4137130, 0.1382410, 0.3730540, 0.3085610, 0.8445550, 0.0764929, 0.2685030, 0.7492750, 0.3044090, 0.5076560, 0.0227180, 0.2494260, 0.1521560, 0.6000770, 0.0236299, 0.0918697, 0.6289560, 0.4593630, 0.4021120, 0.9784450, 0.2027060, 0.3307330, 0.8855350, 0.1042830, 0.3522240, 0.3639500, 0.6031360, 0.1821130, 0.3855590, 0.1451520, 0.4846390, 0.6941100, 0.4597170, 0.4629940, 0.1502520, 0.5867280, 0.9751840, 0.2229700, 0.5277280, 0.1813410, 0.9542980, 0.5175840, 0.3053690, 0.2279530, 0.0774537, 0.0623895, 0.9524640, 0.4914850, 0.4857990, 0.5604000, 0.7049210, 0.9341390, 0.7646320, 0.5200140, 0.4645030, 0.0301845, 0.2824270, 0.0559309, 0.7063850, 0.8377970, 0.6599370, 0.9331040, 0.9453080, 0.2045230, 0.8422190, 0.2267370, 0.9333950, 0.5175320, 0.7578790, 0.9160760, 0.7469880, 0.9229220, 0.4449980, 0.6763780, 0.0094540, 0.2342590, 0.0040166, 0.1486380, 0.0075680, 0.6445940, 0.5203140, 0.3312400, 0.1233810, 0.6449740, 0.0106213, 0.7143200, 0.2191320, 0.8790740, 0.4942060, 0.6439510, 0.9306280, 0.4602340, 0.7181500, 0.5329420, 0.5813610, 0.8621790, 0.8242120, 0.4431260, 0.3833200, 0.8589200, 0.3128730, 0.8365860, 0.2488590, 0.3305430, 0.4424050, 0.6212780, 0.2997030, 0.2796810, 0.9029850, 0.7991840, 0.6486560, 0.7400430, 0.0202659, 0.0571749, 0.3891250, 0.0160444, 0.5603650, 0.2710300, 0.3036670, 0.7713910, 0.6272630, 0.5937740, 0.3796000, 0.1314050, 0.8986940, 0.0346755, 0.5142060, 0.8216660, 0.6680480, 0.8239330, 0.8600900, 0.7700780, 0.2647690, 0.9960680, 0.7752910, 0.2091010, 0.5332120, 0.1010250, 0.5804790, 0.7674280, 0.6884410, 0.9309710, 0.4132980, 0.5911050, 0.6212440, 0.9151900, 0.5417750, 0.6319520, 0.4632780, 0.7969190, 0.4431960, 0.8446090, 0.6569130, 0.9373660, 0.8107010, 0.7748230, 0.4015600, 0.6985390, 0.8261480, 0.9776450, 0.2266680, 0.6831780, 0.0476220, 0.7990130, 0.9653870, 0.8322610, 0.7931950, 0.7705320, 0.6016250, 0.5809500, 0.5744480, 0.6025420, 0.1678080, 0.7808640, 0.0021000, 0.4310650, 0.0202764, 0.4252830, 0.1424460, 0.3484840, 0.2201700, 0.2271960, 0.0519443, 0.0670153, 0.3874240, 0.8885090, 0.8881030, 0.6161330, 0.3263570, 0.4956010, 0.1078270, 0.1359000, 0.0386691, 0.0450091, 0.1359430, 0.6745880, 0.4027270, 0.6942290, 0.6245760, 0.6029850, 0.8521750, 0.6209080, 0.1333660, 0.3557520, 0.2627170, 0.0646071, 0.5407630, 0.0124973, 0.7232120, 0.9532910, 0.7685950, 0.1483780, 0.2077040, 0.4030770, 0.8736990, 0.3684570, 0.2290230, 0.8616150, 0.2267960, 0.6428230, 0.1049960, 0.7701150, 0.5971370, 0.6015390, 0.0061993, 0.4950760, 0.6756710, 0.3660490, 0.9952780, 0.6568520, 0.5795420, 0.9276730, 0.5882040, 0.3427670, 0.5402340, 0.1519320, 0.4874020, 0.9393380, 0.7415860, 0.7102650, 0.8448240, 0.1178210, 0.2857350, 0.8702350, 0.0099742, 0.8071020, 0.3429770, 0.9286890, 0.2840120, 0.3472130, 0.0405582, 0.5633390, 0.1699600, 0.8750190, 0.0279804, 0.6440220, 0.1191350, 0.1444400, 0.0245382, 0.7480850, 0.5016910, 0.5615330, 0.9317580, 0.2913760, 0.3407650, 0.9101610, 0.3564260, 0.7383640, 0.8136830, 0.2868230, 0.4561640, 0.6902130, 0.1840420, 0.4679690, 0.6404870, 0.1957560, 0.2721700, 0.2275550, 0.7170530, 0.8215960, 0.4002780, 0.3780370, 0.1728960, 0.4796630, 0.0877750, 0.7159040, 0.7654720, 0.1411920, 0.2911280, 0.1121760, 0.7815170, 0.0777780, 0.0342828, 0.6245730, 0.1259600, 0.6629980, 0.5919880, 0.3460180, 0.7335800, 0.9477610, 0.8079100, 0.0444241, 0.8715390, 0.7950160, 0.3448870, 0.5739650, 0.6871590, 0.1020760, 0.5260710, 0.3138230, 0.9143850, 0.4996710, 0.1707840, 0.1818680, 0.1439320, 0.4670280, 0.2733560, 0.8116800, 0.3313800, 0.2111440, 0.6671500, 0.8117790, 0.5198900, 0.6790620, 0.3141400, 0.1951690, 0.7294720, 0.7259720, 0.4349700, 0.1108590, 0.1844330, 0.7181340, 0.1094440, 0.2709840, 0.9250700, 0.7569260, 0.9431800, 0.2652650, 0.8857710, 0.9549770, 0.7886410, 0.9084520, 0.3184610, 0.9294640, 0.6758110, 0.9658480, 0.4870440, 0.3840250, 0.4878920, 0.0160075, 0.1265850, 0.0840758, 0.5412280, 0.4356190, 0.2059760, 0.1156660, 0.0103096, 0.5391970, 0.7699970, 0.2482720, 0.5120150, 0.8225120, 0.3600130, 0.2425940, 0.5168880, 0.9987050, 0.9036010, 0.8690720, 0.5166000, 0.6791340, 0.9364790, 0.9219080, 0.0991829, 0.7763010, 0.7309170, 0.5143930, 0.9021310, 0.4349790, 0.7689570, 0.8159200, 0.3394340, 0.1899160, 0.6885280, 0.9235670, 0.2867920, 0.8844140, 0.6476780, 0.6532180, 0.4012660, 0.3219910, 0.3030840, 0.6019840, 0.0600410, 0.7743490, 0.9911680, 0.6051570, 0.3767740, 0.4013380, 0.2222210, 0.4514760, 0.9562650, 0.7572560, 0.8399640, 0.9316500, 0.9114160, 0.0593650, 0.7033740, 0.3911930, 0.7769300, 0.5009410, 0.7506700, 0.5439630, 0.1781090, 0.9061430, 0.0174257, 0.8672990, 0.5254300, 0.1094830, 0.6314700, 0.3939230, 0.4874370, 0.4822290, 0.5335970, 0.4487440, 0.0352250, 0.5891680, 0.9887660, 0.3754300, 0.4365210, 0.8770380, 0.8717270, 0.4104640, 0.2052400, 0.1140760, 0.0953084, 0.3376810, 0.3038450, 0.5767770, 0.4009930, 0.3725630, 0.6179620, 0.1438850, 0.6513020, 0.1508870, 0.0470087, 0.3974610, 0.9766290, 0.7022530, 0.6596390, 0.7840490, 0.5828070, 0.0695546, 0.0811293, 0.0258326, 0.3725470, 0.3215160, 0.6283370, 0.3106610, 0.9849570, 0.3875160, 0.8007740, 0.9571810, 0.4401080, 0.3174350, 0.5846650, 0.7478680, 0.0062299, 0.0579411, 0.1022220, 0.4424290, 0.6233600, 0.3883630, 0.9903260, 0.1396230, 0.2307200, 0.0160327, 0.8287530, 0.5612600, 0.5670550, 0.6091020, 0.4967110, 0.6083740, 0.7601430, 0.2587850, 0.3911380, 0.1899310, 0.0811973, 0.8097900, 0.6658430, 0.2708210, 0.5916970, 0.5305690, 0.5922810, 0.8190990, 0.4018120, 0.1036470, 0.2785020, 0.5497650, 0.0832909, 0.2342630, 0.1744270, 0.8836640, 0.7266790, 0.3421540, 0.6381710, 0.3781130, 0.7428950, 0.9369750, 0.4026680, 0.1945850, 0.9834510, 0.0279463, 0.0707525, 0.9655520, 0.5868360, 0.7511150, 0.3999270, 0.5141220, 0.4091880, 0.6276600, 0.0975324, 0.7867600, 0.0529683, 0.0720765, 0.2010950, 0.8005230, 0.3600280, 0.1488740, 0.4040690, 0.4481550, 0.4439510, 0.1361850, 0.7037450, 0.2960410, 0.2075010, 0.3997570, 0.5355510, 0.9801190, 0.1185160, 0.3544730, 0.3558540, 0.1114660, 0.6801310, 0.6104200, 0.7435930, 0.1838920, 0.3657450, 0.3804120, 0.5644540, 0.7773500, 0.8032880, 0.8206080, 0.2097960, 0.3341130, 0.2940000, 0.9015420, 0.0081535, 0.8905740, 0.9396390, 0.1616070, 0.5218150, 0.7693300, 0.0046586, 0.2654170, 0.6268910, 0.2769680, 0.3057430, 0.8081840, 0.4818340, 0.9930670, 0.4594170, 0.0788334, 0.1619990, 0.6472180, 0.5963010, 0.3409770, 0.9907420, 0.4973450, 0.0538209, 0.1963470, 0.5379350, 0.7206040, 0.4757820, 0.0564678, 0.8359920, 0.7000850, 0.8459170, 0.6310330, 0.3727190, 0.1260880, 0.6525950, 0.4565060, 0.7728110, 0.3250650, 0.1609800, 0.9967960, 0.4248860, 0.8513130, 0.5483310, 0.5641930, 0.0487646, 0.9783770, 0.9943050, 0.0191764, 0.5800090, 0.1644420, 0.9367170, 0.6351340, 0.4587060, 0.0490537, 0.8657760, 0.7223990, 0.7287830, 0.4096380, 0.6447800, 0.2639610, 0.7197410, 0.5238770, 0.4292480, 0.2951760, 0.7541570, 0.0386496, 0.4015090, 0.1969730, 0.1723200, 0.2722920, 0.9137570, 0.2682080, 0.0944083, 0.3398600, 0.3720110, 0.7550490, 0.4028740, 0.2757030, 0.8759390, 0.6679770, 0.6941840, 0.6697170, 0.0323397, 0.9253640, 0.8887650, 0.4101090, 0.9930460, 0.1361780, 0.4457040, 0.8013740, 0.4111790, 0.7054990, 0.9449410, 0.1804920, 0.6636830, 0.9812870, 0.7924080, 0.5968330, 0.3122730, 0.9021120, 0.6773250, 0.8483980, 0.1949160, 0.6193090, 0.8649500, 0.1143260, 0.4601790, 0.4280160, 0.6723250, 0.6378100, 0.1761520, 0.9169270, 0.4712350, 0.8296020, 0.4467770, 0.9246780, 0.4338660, 0.7634010, 0.7477520, 0.5141670, 0.2865240, 0.0674303, 0.4348730, 0.5482950, 0.5616200, 0.1394810, 0.2506930, 0.0792231, 0.6954570, 0.2967850, 0.6185810, 0.1727640, 0.1079510, 0.6691570, 0.1462180, 0.9084860, 0.9073560, 0.1524390, 0.1015940, 0.7526440, 0.0440914, 0.6944870, 0.8206410, 0.2902540, 0.9664710, 0.8320650, 0.3370890, 0.5060190, 0.7383030, 0.1673480, 0.7599160, 0.5982820, 0.8057260, 0.5876320, 0.1255170, 0.4068970, 0.4614890, 0.0546947, 0.0893893, 0.3535940, 0.9268540, 0.0935342, 0.7862810, 0.2585830, 0.4929610, 0.0505512, 0.7359000, 0.2692820, 0.9725290, 0.8130330, 0.9148490, 0.5103490, 0.4526090, 0.2827600, 0.6981670, 0.1923840, 0.4664180, 0.2663510, 0.3333110, 0.0873102, 0.2587710, 0.6352970, 0.6999280, 0.1562920, 0.8272270, 0.3793930, 0.3864410, 0.2127230, 0.5253640, 0.2308400, 0.1768350, 0.1395570, 0.4626540, 0.4677640, 0.6021250, 0.2647550, 0.0432039, 0.6232080, 0.5323690, 0.5362760, 0.9125620, 0.1575890, 0.2018030, 0.6388030, 0.2412790, 0.0935721, 0.9647150, 0.1006100, 0.0151395, 0.1807630, 0.9581900, 0.5021640, 0.2973580, 0.6850120, 0.5680620, 0.9268340, 0.3434440, 0.9217740, 0.2292620, 0.2922360, 0.4061290, 0.4422020, 0.9652240, 0.6557680, 0.9681060, 0.1424770, 0.4704310, 0.8554120, 0.6369300, 0.3425100, 0.3060010, 0.0683669, 0.5944640, 0.0834769, 0.2188230, 0.2694250, 0.0980632, 0.8033720, 0.5066830, 0.4476460, 0.0294077, 0.7180360, 0.5091560, 0.3863140, 0.1214700, 0.3927080, 0.2932910, 0.6284890, 0.4962400, 0.9529960, 0.9173590, 0.3782720, 0.9626610, 0.3520350, 0.1800780, 0.1973760, 0.7248710, 0.3353440, 0.7266170, 0.9951370, 0.3794540, 0.7632550, 0.3016580, 0.6204130, 0.8175660, 0.3257100, 0.5300910, 0.3648150, 0.9225020, 0.6502940, 0.3292770, 0.4483320, 0.2022940, 0.6123560, 0.3689640, 0.0245940, 0.2218170, 0.6291620, 0.5128470, 0.2892840, 0.6108270, 0.6893860, 0.5735930, 0.2014200, 0.3931840, 0.0486366, 0.3986240, 0.7433880, 0.6922420, 0.0499728, 0.6930120, 0.3303580, 0.9247490, 0.8841100, 0.0703700, 0.6288070, 0.8970660, 0.5332270, 0.3091450, 0.2374770, 0.3965410, 0.1859380, 0.5313290, 0.1704160, 0.3465850, 0.5981200, 0.2012750, 0.0681673, 0.3878180, 0.3172690, 0.9839440, 0.9799450, 0.1417040, 0.0099171, 0.9473960, 0.9840760, 0.2777230, 0.0392849, 0.0352798, 0.0943149, 0.9976240, 0.0611254, 0.0391288, 0.7011820, 0.8795180, 0.6973050, 0.3475360, 0.6947180, 0.0254080, 0.0473658, 0.4072930, 0.7044890, 0.5205860, 0.7100460, 0.2679020, 0.6034710, 0.1795280, 0.8876300, 0.2175960, 0.1426860, 0.4477400, 0.3144660, 0.1782390, 0.6623630, 0.4516300, 0.5492990, 0.6181030, 0.3246320, 0.5701350, 0.9636820, 0.9652340, 0.0577224, 0.6083980, 0.4905150, 0.9607970, 0.7008890, 0.5089620, 0.6816150, 0.2367370, 0.5871730, 0.4579290, 0.7153220, 0.3947820, 0.6483250, 0.1229380, 0.7100080, 0.4800800, 0.5151320, 0.3103420, 0.8482150, 0.0115097, 0.7133940, 0.2614500, 0.4008260, 0.2231270, 0.0897239, 0.0094894, 0.8299810, 0.0675502, 0.4172780, 0.2708030, 0.5097350, 0.2474940, 0.9391960, 0.5125170, 0.0235202, 0.8844130, 0.0540106, 0.6745150, 0.5936440, 0.1179910, 0.7889990, 0.4117090, 0.5860720, 0.0853498, 0.7247920, 0.9678720, 0.8628310, 0.3542240, 0.9002370, 0.4046270, 0.2948870, 0.5913430, 0.0607587, 0.4483810, 0.9541920, 0.9814270, 0.6110190, 0.5131570, 0.9183380, 0.0143513, 0.4273990, 0.5001910, 0.0228536, 0.9329900, 0.3340870, 0.2288790, 0.4236030, 0.3115270, 0.5922300, 0.0747541, 0.5989130, 0.6732920, 0.1430020, 0.1833470, 0.1064840, 0.8430170, 0.5797350, 0.3155070, 0.6451030, 0.5664050, 0.9184860, 0.1854750, 0.2125850, 0.9500360, 0.8840290, 0.1619110, 0.6511860, 0.2247230, 0.6644150, 0.2902870, 0.1320890, 0.6977520, 0.4012130, 0.5256570, 0.7584130, 0.3865160, 0.9402190, 0.0019782, 0.5050030, 0.2631490, 0.3850440, 0.9595450, 0.6950050, 0.5415120, 0.1253040, 0.5733380, 0.0845138, 0.9804150, 0.6857450, 0.1985600, 0.7904580, 0.9971510, 0.8235940, 0.9324730, 0.6184770, 0.3232430, 0.6415080, 0.7761480, 0.7207750, 0.7246690, 0.9990340, 0.2724720, 0.1235440, 0.1540990, 0.6916670, 0.7228120, 0.3218540, 0.6365760, 0.2734820, 0.3585550, 0.9914730, 0.8288430, 0.5865600, 0.6681350, 0.4487720, 0.9420290, 0.8122320, 0.9442040, 0.6905970, 0.9219410, 0.9474820, 0.2765560, 0.1809890, 0.6702600, 0.8867870, 0.7803740, 0.7653760, 0.8285700, 0.0597371, 0.6980560, 0.9296280, 0.3703620, 0.2995470, 0.9835380, 0.8901350, 0.1308470, 0.9536370, 0.0619902, 0.6014830, 0.8379440, 0.7190630, 0.2487480, 0.1241330, 0.2603710, 0.5951860, 0.6975130, 0.7016960, 0.7631360, 0.3898470, 0.7319590, 0.9310560, 0.9889760, 0.1258520, 0.9555590, 0.4223190, 0.7638910, 0.2725370, 0.3860450, 0.7589000, 0.2153160, 0.1335290, 0.4254760, 0.7987810, 0.6640640, 0.7647820, 0.0015695, 0.9057530, 0.4736930, 0.3972490, 0.8668450, 0.7828120, 0.3726150, 0.7891530, 0.2566250, 0.5296370, 0.0610593, 0.4443960, 0.1512180, 0.2462730, 0.9915970, 0.1090550, 0.5283070, 0.5068540, 0.0562730, 0.9824450, 0.6897040, 0.8177550, 0.5943070, 0.5580590, 0.6899610, 0.9541940, 0.6938890, 0.8858770, 0.1965490, 0.1321620, 0.4941940, 0.8370090, 0.2533520, 0.4695890, 0.9374020, 0.5060690, 0.3550800, 0.1501900, 0.6746690, 0.6862980, 0.7163260, 0.9192100, 0.9026580, 0.7726290, 0.2742970, 0.6578880, 0.2575500, 0.2605210, 0.0536524, 0.9747520, 0.8189380, 0.8512580, 0.9693230, 0.8496760, 0.1084130, 0.6433380, 0.3389490, 0.7581810, 0.2526000, 0.4821550, 0.1751500, 0.3119460, 0.9038050, 0.4294420, 0.9665870, 0.9408750, 0.3523780, 0.2090970, 0.5009810, 0.2864980, 0.7493820, 0.2950710, 0.5543530, 0.7601390, 0.9385800, 0.2652270, 0.9942620, 0.1471980, 0.5878890, 0.5441030, 0.7895980, 0.2410650, 0.7209760, 0.9033380, 0.8547790, 0.5828550, 0.6810760, 0.4335560, 0.7923370, 0.2144880, 0.5433650, 0.2237820, 0.2470670, 0.4658720, 0.0756143, 0.4012210, 0.5670660, 0.5502220, 0.1081130, 0.1514850, 0.6065610, 0.7238760, 0.1114270, 0.7785880, 0.7681590, 0.1499110, 0.0059389, 0.2630620, 0.9967180, 0.8207220, 0.0999561, 0.7656770, 0.3949100, 0.6871100, 0.7437380, 0.5144240, 0.8344960, 0.3059900, 0.1060730, 0.1088490, 0.1637970, 0.2663330, 0.3051170, 0.2009190, 0.1945110, 0.7667110, 0.6550970, 0.1552670, 0.5135020, 0.5022780, 0.9979660, 0.1732610, 0.4610580, 0.5316570, 0.9417340, 0.7801650, 0.4042490, 0.7878990, 0.0331769, 0.9438240, 0.6906600, 0.3363680, 0.0709532, 0.3468950, 0.7838490, 0.0021231, 0.3406110, 0.0268374, 0.8030730, 0.4337860, 0.2373690, 0.8551890, 0.0025808, 0.6639180, 0.8748950, 0.2093230, 0.9261020, 0.6114200, 0.0697385, 0.8821280, 0.9657740, 0.3730850, 0.3014390, 0.1283160, 0.4752300, 0.1635610, 0.9838330, 0.6431800, 0.9863560, 0.7228600, 0.2970090, 0.1037600, 0.3138450, 0.7882810, 0.7507470, 0.2235520, 0.1994370, 0.5732010, 0.5472950, 0.1523960, 0.2213770, 0.8936120, 0.0168712, 0.3288280, 0.2211280, 0.6751350, 0.5519800, 0.4526020, 0.4179590, 0.0040056, 0.4670670, 0.1303090, 0.8155870, 0.1118400, 0.8991280, 0.1368980, 0.6428140, 0.5909770, 0.4997330, 0.3682430, 0.1137550, 0.0959078, 0.0692972, 0.5941720, 0.3352730, 0.6888380, 0.3568610, 0.3329040, 0.6609200, 0.1117310, 0.3756910, 0.5606760, 0.4012910, 0.2984950, 0.5799880, 0.5776480, 0.6486580, 0.8936940, 0.1841640, 0.5297140, 0.8741020, 0.2013400, 0.2713440, 0.0011868, 0.7137630, 0.8521240, 0.8041440, 0.1169840, 0.3849810, 0.7189480, 0.7326120, 0.9566820, 0.2989380, 0.3062740, 0.5168990, 0.8849890, 0.8976650, 0.4962450, 0.3769900, 0.0233866, 0.1739690, 0.6783090, 0.8666600, 0.0822737, 0.7554740, 0.5892600, 0.2151310, 0.8617170, 0.7531930, 0.6468350, 0.0594414, 0.1059990, 0.9081290, 0.6232850, 0.3350880, 0.4984580, 0.3487300, 0.8770410, 0.4664800, 0.2392150, 0.0375377, 0.8793530, 0.7374710, 0.5278570, 0.3899630, 0.7294870, 0.5055200, 0.9987860, 0.5090390, 0.4058960, 0.5095730, 0.1773760, 0.1864990, 0.2127110, 0.3384130, 0.0186218, 0.5788500, 0.0395564, 0.2169370, 0.4108910, 0.2662530, 0.2934810, 0.7606650, 0.1156990, 0.4427970, 0.4885540, 0.9541000, 0.3851010, 0.2585500, 0.0604153, 0.0924547, 0.2332740, 0.3486330, 0.6283100, 0.2855750, 0.8083950, 0.5611440, 0.5024140, 0.9558770, 0.6857060, 0.7549880, 0.4075650, 0.6374560, 0.6384980, 0.4894190, 0.7382240, 0.2251570, 0.9101300, 0.0373303, 0.0671782, 0.2925690, 0.8477730, 0.9955480, 0.0188255, 0.5613020, 0.3736500, 0.1304100, 0.2289210, 0.3343480, 0.7265210, 0.5270450, 0.0207100, 0.6253360, 0.1072220, 0.3420270, 0.3120370, 0.5339230, 0.8525590, 0.3710180, 0.1522940, 0.1738170, 0.9856940, 0.9909300, 0.4252230, 0.6310430, 0.0708148, 0.4448940, 0.8264210, 0.7688160, 0.2342140, 0.3905100, 0.7830270, 0.3199690, 0.2655050, 0.2264060, 0.9553160, 0.1948030, 0.0345524, 0.6072520, 0.1816020, 0.8838550, 0.2996590, 0.2967710, 0.2748080, 0.3924660, 0.0226123, 0.8360040, 0.5845130, 0.4805100, 0.9839280, 0.9949630, 0.2586500, 0.9883280, 0.9188970, 0.7277180, 0.5934600, 0.1981100, 0.1255590, 0.8762200, 0.1427400, 0.0923326, 0.3029980, 0.5771690, 0.5806870, 0.0260272, 0.5179030, 0.8915560, 0.1248840, 0.3133100, 0.2814550, 0.6081440, 0.8693970, 0.4187220, 0.2698480, 0.8948010, 0.9389350, 0.2543970, 0.9099630, 0.9100800, 0.9657490, 0.9978740, 0.2492640, 0.7749230, 0.2266600, 0.3361180, 0.1780730, 0.6981950, 0.3189340, 0.4854910, 0.6524080, 0.0281007, 0.1885550, 0.8255900, 0.9316340, 0.5602800, 0.9029590, 0.5246330, 0.3887920, 0.7092010, 0.1811620, 0.4524370, 0.4962900, 0.1564060, 0.8295370, 0.0594514, 0.0661466, 0.4066640, 0.6977710, 0.3564360, 0.5263990, 0.9847150, 0.8461340, 0.6224430, 0.3112100, 0.2814500, 0.1984650, 0.5467730, 0.3826040, 0.0237089, 0.7431600, 0.0896665, 0.6653870, 0.1767840, 0.9433970, 0.1921440, 0.3878050, 0.1430450, 0.5377090, 0.7373430, 0.2629910, 0.4085910, 0.5753620, 0.6573880, 0.6243580, 0.9472190, 0.6310810, 0.7329550, 0.3960680, 0.0072950, 0.6746710, 0.2142820, 0.3874810, 0.3366010, 0.1085510, 0.5217040, 0.7612800, 0.6268970, 0.3571330, 0.6220930, 0.3281020, 0.3127150, 0.4716210, 0.2406920, 0.6294350, 0.3764380, 0.9024370, 0.9044030, 0.3864810, 0.4574290, 0.9248130, 0.5140700, 0.4851120, 0.7409150, 0.3131900, 0.7756240, 0.7465640, 0.6418780, 0.5924490, 0.4224650, 0.3373970, 0.7890890, 0.7414770, 0.8899260, 0.6205810, 0.7715480, 0.2007730, 0.0224243, 0.6278590, 0.5090430, 0.8647530, 0.5879950, 0.1219100, 0.5784320, 0.5450500, 0.6640110, 0.2692960, 0.0144626, 0.6056110, 0.2947460, 0.0718636, 0.3305410, 0.0499776, 0.1411190, 0.2882690, 0.2410710, 0.4400780, 0.7953110, 0.7101640, 0.5566740, 0.4890210, 0.0367743, 0.2479610, 0.0747430, 0.6109450, 0.1588980, 0.2418870, 0.1714300, 0.8592690, 0.5592470, 0.8150700, 0.8204730, 0.2702690, 0.9564510, 0.1567270, 0.6111830, 0.9433950, 0.7830260, 0.3080010, 0.7807270, 0.7554470, 0.2663120, 0.5553010, 0.2429540, 0.5447430, 0.3687010, 0.1531340, 0.1047130, 0.7453280, 0.5124190, 0.3241720, 0.4353590, 0.2211670, 0.3775170, 0.9916820, 0.1620050, 0.7116460, 0.4297190, 0.3230200, 0.3569010, 0.0390569, 0.2744480, 0.4480660, 0.9098220, 0.1287040, 0.7298730, 0.3694950, 0.8581680, 0.3285810, 0.6453340, 0.8138680, 0.3126460, 0.1893730, 0.4234730, 0.1061980, 0.1828110, 0.0744468, 0.3475120, 0.8881380, 0.6503170, 0.9405250, 0.8202320, 0.1937450, 0.4597900, 0.0928449, 0.5723780, 0.6572270, 0.6196420, 0.8193340, 0.8721010, 0.3675210, 0.5975880, 0.8469860, 0.0881379, 0.7356970, 0.9469610, 0.0668435, 0.9510170, 0.5632600, 0.8441910, 0.0051679, 0.8413210, 0.1944340, 0.5760520, 0.3278480, 0.4151400, 0.8104830, 0.1702260, 0.5006220, 0.8415750, 0.8550480, 0.0836501, 0.4746020, 0.1579540, 0.3317340, 0.1817210, 0.2649720, 0.0646802, 0.1244630, 0.3847370, 0.0067872, 0.5895460, 0.8055080, 0.7826130, 0.2013730, 0.5635350, 0.2325570, 0.5881820, 0.0998175, 0.2283320, 0.6095520, 0.7946270, 0.4423650, 0.0336123, 0.1274130, 0.9943250, 0.7288430, 0.1056540, 0.0931000, 0.2216070, 0.4693430, 0.6233060, 0.3880930, 0.6500330, 0.5146820, 0.3216340, 0.3530970, 0.4511740, 0.7347270, 0.9870220, 0.7286780, 0.9407670, 0.9029230, 0.4128020, 0.4928480, 0.0117259, 0.5158110, 0.9319450, 0.4534930, 0.9037510, 0.0653333, 0.3440930, 0.4411360, 0.4346250, 0.8741540, 0.6308510, 0.8786790, 0.1764270, 0.8946940, 0.7381230, 0.8997440, 0.9564830, 0.9038440, 0.7733660, 0.4502270, 0.1455900, 0.9851600, 0.1646910, 0.0031155, 0.1696680, 0.1941350, 0.0192863, 0.3532120, 0.1321330, 0.4303470, 0.4970510, 0.2430670, 0.2177900, 0.3740440, 0.1629570, 0.2499810, 0.8667330, 0.0705503, 0.0027678, 0.0354401, 0.6207550, 0.5467060, 0.6422110, 0.4687960, 0.2162460, 0.1524840, 0.0857022, 0.6267270, 0.4590980, 0.7320680, 0.9346080, 0.8328770, 0.2522410, 0.3535130, 0.4847060, 0.4363190, 0.5519930, 0.7500680, 0.1616170, 0.3431100, 0.1981380, 0.8950640, 0.4764970, 0.7383730, 0.8198900, 0.1436160, 0.6459620, 0.4276260, 0.5180440, 0.7660530, 0.4925970, 0.9354560, 0.7012280, 0.0850516, 0.1477460, 0.2548520, 0.0077067, 0.4998510, 0.5684250, 0.5586210, 0.9227440, 0.7139860, 0.4787920, 0.2675560, 0.2775030, 0.6904630, 0.4975710, 0.6635750, 0.7914070, 0.4424440, 0.5400100, 0.2628160, 0.0344078, 0.7751210, 0.9847490, 0.5114180, 0.8968250, 0.1516410, 0.2228920, 0.5624620, 0.0418695, 0.1130320, 0.0046975, 0.8447880, 0.0048562, 0.5960620, 0.4313710, 0.6853910, 0.8488930, 0.9530650, 0.6633300, 0.3247750, 0.0482924, 0.9411870, 0.2438960, 0.8511580, 0.3679400, 0.0968893, 0.7731470, 0.7483640, 0.5633240, 0.8877430, 0.2897910, 0.6387570, 0.6698470, 0.1338030, 0.8311510, 0.6348650, 0.6206600, 0.6441150, 0.9225490, 0.8297640, 0.9443350, 0.0492086, 0.0598250, 0.1146800, 0.8663100, 0.7550870, 0.1124790, 0.5905840, 0.8867160, 0.1631950, 0.9178910, 0.2702930, 0.2468280, 0.0461997, 0.8212920, 0.3839270, 0.5922680, 0.5909710, 0.9854710, 0.8658860, 0.1078680, 0.3163630, 0.6863420, 0.6708680, 0.0355104, 0.5879850, 0.3204140, 0.5822750, 0.8054990, 0.1901980, 0.3750820, 0.1705350, 0.1395890, 0.0920875, 0.3687330, 0.2242380, 0.9023150, 0.9877700, 0.1059010, 0.2169810, 0.9012520, 0.0154705, 0.2781610, 0.0467885, 0.0197655, 0.4963860, 0.1490130, 0.5998810, 0.4424520, 0.2247180, 0.0092350, 0.8775790, 0.7509590, 0.5634700, 0.9533570, 0.9052740, 0.5749590, 0.8782240, 0.6161180, 0.7047450, 0.2094630, 0.6244000, 0.2583050, 0.3182590, 0.9670720, 0.3086500, 0.7611730, 0.8978890, 0.7963160, 0.6873890, 0.7602140, 0.6411920, 0.4272750, 0.3065350, 0.3832750, 0.4601360, 0.0953929, 0.6330440, 0.5152900, 0.1779940, 0.1846950, 0.6620860, 0.6886720, 0.8532580, 0.2272490, 0.1068230, 0.6582580, 0.0897870, 0.4923490, 0.9047110, 0.0051937, 0.6762720, 0.4101160, 0.9435750, 0.8753460, 0.4793050, 0.3879890, 0.6072320, 0.3859910, 0.4748990, 0.3746120, 0.8730050, 0.1783370, 0.5281440, 0.5350820, 0.9731060, 0.5446980, 0.3157400, 0.2592250, 0.2890660, 0.3599570, 0.8503720, 0.7631550, 0.0810297, 0.2968880, 0.5231600, 0.4481580, 0.1942020, 0.8530370, 0.7114600, 0.4988370, 0.3351890, 0.3357620, 0.7523330, 0.0745497, 0.9790390, 0.4933010, 0.7873570, 0.5317550, 0.1608920, 0.2956830, 0.2830060, 0.9040950, 0.3330890, 0.2492080, 0.3569710, 0.2234840, 0.7720440, 0.4169650, 0.5832730, 0.4731490, 0.2103330, 0.7193440, 0.1664530, 0.1346010, 0.3917440, 0.6398030, 0.8521720, 0.4628410, 0.1041940, 0.4633620, 0.7696810, 0.2891010, 0.9646030, 0.4363480, 0.0876910, 0.6224150, 0.2415180, 0.0057658, 0.2242650, 0.6456620, 0.8128750, 0.2804420, 0.1940670, 0.0127567, 0.7947130, 0.7267310, 0.4228260, 0.9979530, 0.0699841, 0.2532890, 0.1592940, 0.0899736, 0.6422130, 0.2585520, 0.2763750, 0.8357830, 0.1335810, 0.6391710, 0.2024160, 0.4593320, 0.7546290, 0.3540040, 0.0676632, 0.8409670, 0.3156530, 0.7813270, 0.8189590, 0.9775050, 0.0556196, 0.7371110, 0.4445510, 0.4867060, 0.6835660, 0.7284170, 0.0068706, 0.2279430, 0.1692620, 0.7170460, 0.8259380, 0.3420010, 0.7497990, 0.7991860, 0.4831920, 0.1735390, 0.4537990, 0.3265880, 0.1211680, 0.2965230, 0.7874410, 0.0669131, 0.1021410, 0.3091770, 0.2477700, 0.8527590, 0.4247480, 0.5653140, 0.2242000, 0.6363470, 0.1979850, 0.3676470, 0.5525700, 0.2898320, 0.9194250, 0.6193910, 0.3758970, 0.8113510, 0.7843390, 0.9150010, 0.0819345, 0.2608680, 0.0724862, 0.7906520, 0.0146286, 0.8898050, 0.3849050, 0.0999590, 0.4756150, 0.2254880, 0.2158640, 0.0013373, 0.2449740, 0.8493100, 0.1919980, 0.0865416, 0.8002820, 0.4473960, 0.0349332, 0.5748180, 0.4177360, 0.9855740, 0.5345390, 0.7039820, 0.6481140, 0.3249930, 0.3828090, 0.1601250, 0.5144310, 0.5226810, 0.7392030, 0.9913150, 0.9186170, 0.8812290, 0.8562620, 0.0344090, 0.5299830, 0.8423540, 0.9246350, 0.0745926, 0.9175070, 0.2316900, 0.8081040, 0.5868900, 0.8750580, 0.6326160, 0.0123006, 0.4631190, 0.1652820, 0.0411444, 0.1412320, 0.2440110, 0.4951630, 0.1573670, 0.9724490, 0.2758710, 0.6532560, 0.0684292, 0.6610630, 0.5959930, 0.7477160, 0.7436860, 0.5146670, 0.8282460, 0.2047110, 0.3026700, 0.4440070, 0.0519424, 0.2982110, 0.3707150, 0.0164968, 0.8084940, 0.7616030, 0.2817020, 0.3699820, 0.6940910, 0.0393768, 0.1915540, 0.9293910, 0.2812620, 0.9839630, 0.2840670, 0.5040720, 0.1168300, 0.3829590, 0.9129470, 0.7211830, 0.5717790, 0.8271240, 0.3571970, 0.9893070, 0.2854670, 0.3913660, 0.1203400, 0.7963540, 0.1499640, 0.2343730, 0.7371340, 0.8102780, 0.3624880, 0.9300510, 0.1318330, 0.1972740, 0.4972180, 0.0854875, 0.0956049, 0.5711640, 0.0547849, 0.2758760, 0.5001440, 0.2989470, 0.6812780, 0.4386600, 0.9523000, 0.8111450, 0.6782420, 0.4743620, 0.2521000, 0.0822533, 0.1033280, 0.6504920, 0.8639670, 0.0001646, 0.1048860, 0.8706430, 0.4598670, 0.7703220, 0.3723100, 0.7356540, 0.0357558, 0.9936870, 0.1072880, 0.3902270, 0.1771350, 0.3741170, 0.1509670, 0.1319940, 0.6264530, 0.6154480, 0.3556980, 0.3544270, 0.2280310, 0.0086045, 0.2990430, 0.0516253, 0.4432200, 0.6602410, 0.1638160, 0.1391590, 0.6151970, 0.3956990, 0.0843927, 0.7229610, 0.4813430, 0.9468080, 0.9117370, 0.0194119, 0.5611690, 0.2866660, 0.0326114, 0.3202930, 0.3047980, 0.2833830, 0.7407690, 0.6776100, 0.7382690, 0.8835430, 0.1363110, 0.0643888, 0.9309500, 0.0234121, 0.4336830, 0.9154960, 0.1142520, 0.1966400, 0.2152250, 0.4392960, 0.9470380, 0.6262830, 0.8377920, 0.3593160, 0.5154830, 0.9033030, 0.7841330, 0.2861750, 0.2645370, 0.8416070, 0.1173600, 0.9769400, 0.7871540, 0.0430673, 0.2346290, 0.6233080, 0.2287270, 0.9345000, 0.3965720, 0.1522510, 0.8885020, 0.7341700, 0.1418020, 0.2924590, 0.8793740, 0.6063140, 0.7410150, 0.5315020, 0.5155460, 0.7625500, 0.6359050, 0.7623200, 0.5718010, 0.4303810, 0.1188080, 0.8490030, 0.9818700, 0.5888760, 0.3023120, 0.0950337, 0.7545320, 0.3911800, 0.5577450, 0.6701150, 0.6029400, 0.9652090, 0.5405540, 0.7124950, 0.2537520, 0.5967210, 0.4162570, 0.5273840, 0.8331670, 0.0464175, 0.0989103, 0.6669570, 0.2747010, 0.6972900, 0.0587434, 0.9782650, 0.9965620, 0.4407890, 0.4519890, 0.5629660, 0.2955860, 0.8357000, 0.4209090, 0.4978350, 0.2061670, 0.4361330, 0.6912480, 0.3560640, 0.6937410, 0.5118960, 0.7244010, 0.5430630, 0.3212620, 0.9121490, 0.7361140, 0.7807190, 0.4367510, 0.5613460, 0.4140270, 0.7057840, 0.0371946, 0.2403880, 0.9231870, 0.7127470, 0.7680580, 0.3828300, 0.1641800, 0.2830810, 0.5710970, 0.4300000, 0.0627110, 0.6209070, 0.5036890, 0.0077011, 0.4523210, 0.0029354, 0.2151600, 0.1060240, 0.9373460, 0.7607010, 0.7247800, 0.2087200, 0.4005850, 0.3378640, 0.5349830, 0.2833120, 0.1938950, 0.2785860, 0.9385400, 0.6003060, 0.9951260, 0.9239020, 0.1597880, 0.8991380, 0.5956720, 0.3476410, 0.0059898, 0.1885460, 0.6217270, 0.5414400, 0.6117280, 0.7740560, 0.0899378, 0.9196150, 0.6629460, 0.7550210, 0.9673900, 0.5753760, 0.3448740, 0.2854240, 0.8880670, 0.7433620, 0.0932783, 0.0830703, 0.8386430, 0.5207910, 0.5399290, 0.3911440, 0.4775630, 0.7143900, 0.8530210, 0.8255710, 0.7702860, 0.6936570, 0.9508410, 0.2925610, 0.7605690, 0.1170520, 0.1699550, 0.0272872, 0.9401800, 0.4870220, 0.3719700, 0.5925280, 0.4383840, 0.5538310, 0.9703260, 0.9346940, 0.3251220, 0.3770310, 0.1164470, 0.9277290, 0.8386170, 0.6754820, 0.3794290, 0.3352000, 0.6335750, 0.9725530, 0.8639060, 0.9513870, 0.4315320, 0.0701333, 0.9135840, 0.2557460, 0.6727200, 0.9895930, 0.9637080, 0.4160600, 0.2468050, 0.9146060, 0.8212470, 0.0434056, 0.7036910, 0.4572880, 0.3129530, 0.1061150, 0.3862520))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s49,
    done => done_s50,
    start => start_s51,
    ack => ack_s52,
    in_a => in_a_s53,
    out_a => out_a_s54,
    out_offset => out_offset_s55,
    simd_offset => simd_offset_s56,
    op_argument => op_argument_s57,
    op_result => op_result_s58,
    op_send => op_send_s59,
    op_receive => op_receive_s60
);
conv_to_fc_interlayer_u114 : conv_to_fc_interlayer generic map(
    channels => 10,
    channel_width => 8,
    layer_size => 7,
    fc_simd => 10
) port map(
    clk => clk,
    ready => ready_s115,
    done => done_s116,
    start => start_s117,
    ack => ack_s118,
    din => din_s119,
    dout => dout_s120,
    wr_addr => wr_addr_s121,
    rd_addr => rd_addr_s122,
    wren_in => wren_in_s123
);
bias_op_u61 : bias_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 13, frac => 15)),
    bias_spec => fixed_spec(fixed_spec'(int => 1, frac => 11)),
    biases => reals(reals'( 0.9110350, 0.6515300, 0.2094400, 0.0287224, 0.3006430, 0.1099270, 0.6336950, 0.1806030, 0.3290790, 0.2056470))
) port map(
    input => input_s62,
    offset => offset_s63,
    output => output_s64,
    op_send => op_send_s65,
    op_receive => op_receive_s66
);
sigmoid_op_u67 : sigmoid_op generic map(
    input_spec => fixed_spec(fixed_spec'(int => 14, frac => 15)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    step_precision => 2,
    bit_precision => 16
) port map(
    clk => clk,
    input => input_s68,
    output => output_s69,
    op_send => op_send_s70,
    op_receive => op_receive_s71
);

din_s87 <= dout_s7;
ack_s4 <= load_done_s17;
done_s85 <= done_s2;
ready_s74 <= ready_s1;
rd_addr_s80 <= addr_s8;
start_s3 <= start_s76;
din_s6 <= dout_s78;
row_s91 <= row_s10;
wren_s92 <= wren_s11;
wr_addr_s89 <= out_addr_s9;
din_s97 <= dout_s19;
ack_s16 <= load_done_s29;
done_s95 <= done_s14;
ready_s84 <= ready_s13;
rd_addr_s90 <= addr_s20;
start_s15 <= start_s86;
din_s18 <= dout_s88;
row_s101 <= row_s22;
wren_s102 <= wren_s23;
wr_addr_s99 <= out_addr_s21;
din_s107 <= dout_s31;
ack_s28 <= load_done_s41;
done_s105 <= done_s26;
ready_s94 <= ready_s25;
rd_addr_s100 <= addr_s32;
start_s27 <= start_s96;
din_s30 <= dout_s98;
row_s111 <= row_s34;
wren_s112 <= wren_s35;
wr_addr_s109 <= out_addr_s33;
din_s119 <= dout_s43;
ack_s40 <= ack_s118;
done_s116 <= done_s38;
ready_s104 <= ready_s37;
rd_addr_s110 <= addr_s44;
start_s39 <= start_s106;
din_s42 <= dout_s108;
wren_in_s123 <= wren_s47;
wr_addr_s121 <= out_addr_s45;
in_a_s53 <= dout_s120;
start_s51 <= start_s117;
ready_s115 <= ready_s49;
rd_addr_s122 <= std_logic_vector(resize(unsigned(simd_offset_s56), rd_addr_s122'length));
input_s62 <= op_argument_s57;
op_receive_s66 <= op_send_s59;
op_receive_s60 <= op_send_s70;
input_s68 <= output_s64;
op_receive_s71 <= op_send_s65;
offset_s63 <= out_offset_s55;
op_result_s58 <= resize(output_s69, mk(fixed_spec(fixed_spec'(int => 2, frac => 8))));

uPS : ps_clk port map(
    clk => clk,
    rst => rst_sink
);
done_s75 <= start;
test_out <= shift_range(std_logic_vector(get(out_a_s54, to_integer(sel), mk(fixed_spec(fixed_spec'(int => 2, frac => 8))))), 8)(test_out'range) when to_integer(sel) < 10 else "00000000";
end system;
