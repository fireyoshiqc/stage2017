use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library ieee_proposed;
use ieee_proposed.fixed_pkg.all;

library work;
use work.util.all;

entity system is
port(
    start : in std_logic;
    test_out : out std_logic_vector(8 - 1 downto 0);
    sel : in unsigned(8 - 1 downto 0)
);
end system;

architecture system of system is

component fc_layer is
generic(
    input_width : integer;
    output_width : integer;
    simd_width : integer;
    input_spec : fixed_spec;
    weight_spec : fixed_spec;
    op_arg_spec : fixed_spec;
    output_spec : fixed_spec;
    n_weights : integer;
    weights_filename : string;
    weight_values : reals
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : out std_logic;
    done : out std_logic;
    start : in std_logic;
    ack : in std_logic;
    in_a : in std_logic_vector;
    out_a : out std_logic_vector;
    out_offset : out unsigned;
    op_argument : out sfixed;
    op_result : in sfixed;
    op_send : out std_logic;
    op_receive : in std_logic
);
end component;

component interlayer is
generic(
    width : integer;
    word_size : integer
);
port(
    clk : in std_logic;
    rst : in std_logic;
    ready : in std_logic;
    done : in std_logic;
    start : out std_logic;
    ack : out std_logic;
    previous_a : in std_logic_vector;
    next_a : out std_logic_vector
);
end component;




signal ready_s1 : std_logic;
signal done_s2 : std_logic;
signal start_s3 : std_logic;
signal ack_s4 : std_logic;
signal in_a_s5 : std_logic_vector(503 downto 0);
signal out_a_s6 : std_logic_vector(399 downto 0);
signal out_offset_s7 : unsigned(5 downto 0);
signal op_argument_s8 : sfixed(10 downto -14);
signal op_result_s9 : sfixed(1 downto -8);
signal op_send_s10 : std_logic;
signal op_receive_s11 : std_logic;



signal ready_s14 : std_logic;
signal done_s15 : std_logic;
signal start_s16 : std_logic;
signal ack_s17 : std_logic;
signal previous_a_s18 : std_logic_vector(503 downto 0);
signal next_a_s19 : std_logic_vector(503 downto 0);


component ps is
port(
    clk, rst : out std_logic
);
end component;

signal clk, rst_sink : std_logic;
constant rst : std_logic := '0';

function to_vec(r : reals) return std_logic_vector is
    constant input_spec : fixed_spec := fixed_spec(fixed_spec'(int => 1, frac => 8));
    variable ret : std_logic_vector(56 * size(input_spec) - 1 downto 0);
begin
    for i in r'range loop
        ret((1 + i) * size(input_spec) - 1 downto i * size(input_spec)) :=
            std_logic_vector(to_sfixed(r(i), mk(input_spec)));
    end loop;
    return ret;
end to_vec;

begin

fc_layer_u0 : fc_layer generic map(
    input_width => 56,
    output_width => 40,
    simd_width => 14,
    input_spec => fixed_spec(fixed_spec'(int => 1, frac => 8)),
    weight_spec => fixed_spec(fixed_spec'(int => 2, frac => 6)),
    op_arg_spec => fixed_spec(fixed_spec'(int => 11, frac => 14)),
    output_spec => fixed_spec(fixed_spec'(int => 2, frac => 8)),
    n_weights => 2240,
    weights_filename => "whatever",
    weight_values => reals(reals'( 0.0000408, 0.0001156, -0.0007705, -0.0003351, -0.0000950, -0.0000820, 0.0004032, 0.0004182, 0.0003001, -0.0001907, 0.0000297, 0.0001292, 0.0016181, 0.0033509, -0.0004116, 0.0003559, -0.0004802, 0.0006479, 0.0000861, 0.0001580, -0.0002336, -0.0007931, 0.0001428, 0.0002428, 0.0001890, 0.0001554, 0.0000769, -0.0002156, -0.0003911, 0.0005581, -0.0002465, 0.0002428, -0.0002677, 0.0001292, 0.0038330, 0.0061119, 0.0063058, 0.0006660, 0.0018109, 0.0006858, 0.0013706, -0.0008381, -0.0072303, -0.0185001, -0.0347154, -0.0061202, 0.0011924, 0.0005082, 0.0053583, 0.0091062, 0.0035945, 0.0034690, -0.0000003, -0.0001222, -0.0000568, 0.0004877, -0.0001252, 0.0003127, -0.0004140, -0.0001421, -0.0000033, 0.0006630, 0.0109417, 0.0252189, 0.0151279, 0.0068338, 0.0396617, 0.0650002, 0.0643596, 0.0811151, 0.0860193, -0.0110326, -0.0857354, -0.0706970, -0.0742991, -0.0005925, 0.0023063, 0.0138023, 0.0146258, 0.0043074, 0.0012573, -0.0001469, 0.0000623, 0.0000403, -0.0004547, -0.0000152, -0.0005816, -0.0001612, -0.0031084, 0.0046655, 0.0184095, 0.0547722, 0.0458653, 0.0764468, 0.0815437, 0.1466200, 0.0937492, 0.0375963, 0.0035690, -0.1021800, -0.2487210, -0.3082000, -0.2899820, -0.0337810, 0.0001316, 0.0216308, 0.0618042, 0.0580215, 0.0566176, 0.0078293, 0.0029489, 0.0002086, 0.0003119, 0.0001715, -0.0005010, -0.0004678, 0.0152223, 0.0533587, 0.0362833, 0.0299187, 0.0700633, 0.0895389, 0.1649460, 0.1331820, 0.1819780, 0.0565010, -0.1609890, -0.4032590, -0.4190330, -0.3572230, -0.1928310, 0.0605936, 0.0882286, 0.0867366, 0.1055950, 0.0875757, -0.0268386, -0.0430774, -0.0172364, 0.0036921, 0.0001532, 0.0001673, -0.0000059, -0.0072398, 0.0208059, 0.1688750, 0.1909760, 0.0865629, 0.1039180, 0.2798850, 0.3238080, 0.1378940, 0.2829040, -0.2263370, -0.6018320, -0.8534070, -0.5163420, -0.0100411, 0.1574760, 0.2480940, 0.0461678, 0.0378534, 0.0724771, 0.1342370, 0.0580798, -0.0394766, 0.0024487, 0.0076129, 0.0000928, 0.0003728, -0.0064206, -0.0605344, -0.0266544, 0.1227010, 0.1451860, 0.1449620, 0.2019420, 0.2780500, 0.1807230, 0.2340500, 0.1263620, -0.1964740, -0.9113080, -1.1540300, -0.4700730, 0.0665744, 0.1417590, 0.2358060, 0.1873120, -0.0416665, 0.0090010, 0.1549920, 0.0240485, -0.0267736, 0.0006723, 0.0077243, -0.0000285, 0.0023462, -0.0025640, -0.0657071, -0.0152877, 0.0693240, 0.0630817, 0.0741730, 0.0615562, 0.2631320, 0.3346370, 0.2321780, -0.0041563, -0.3724530, -0.8663880, -0.8247520, -0.2379330, 0.0877544, 0.1769310, 0.2037680, 0.1364920, 0.0265569, 0.0691599, 0.0900181, -0.1163740, -0.0665033, 0.0174623, 0.0040099, 0.0009015, 0.0038694, 0.0061569, -0.0065498, 0.0100425, 0.0665915, 0.0086675, 0.1650280, 0.1150910, 0.2559440, 0.2103880, 0.3606190, 0.3568610, -0.2033450, -0.8553220, -0.5303120, 0.0843481, 0.2036230, 0.1661590, 0.1818670, -0.0499374, -0.0155624, -0.0014863, -0.0768179, -0.1490330, -0.0253135, -0.0357896, -0.0058015, -0.0002553, 0.0029923, 0.0110067, 0.0237443, 0.0846660, 0.0344682, -0.0391484, 0.0321596, 0.2034950, 0.0690879, 0.0916413, 0.3515740, 0.4030360, -0.3933870, -0.8713900, -0.0857388, 0.3325590, 0.2552340, 0.1656670, 0.1179140, 0.0361244, 0.0444135, 0.0276070, -0.0936895, -0.0007871, -0.0660689, -0.0471792, 0.0069456, 0.0001135, 0.0033795, 0.0222199, 0.0046883, 0.1319100, 0.0727055, -0.2025440, -0.0965611, 0.1306940, 0.0372889, 0.0024322, 0.3224870, 0.1386070, -0.7207660, -0.6768400, -0.0494575, 0.2243560, 0.2467750, 0.0564180, 0.1677640, -0.0048336, 0.1933900, 0.0008101, -0.0728858, 0.0831703, 0.0314235, -0.0194856, -0.0025027, 0.0003479, 0.0041175, 0.0050364, -0.0131561, 0.0649843, 0.0597026, -0.1620470, -0.2529410, -0.1225150, -0.2856400, -0.1759120, -0.0267279, -0.1076350, -0.4435970, -0.0710733, -0.0131802, 0.1068500, 0.0843650, 0.1885230, -0.0146504, -0.0342709, 0.1375340, -0.0521685, -0.0173079, 0.0171801, 0.0077618, -0.0231124, -0.0034051, 0.0001255, 0.0022242, 0.0204442, -0.0053252, 0.0119030, -0.0699116, -0.0808024, -0.0198391, -0.0490748, -0.3275890, -0.0885521, -0.0497274, -0.2151700, -0.2163290, -0.0213713, 0.1578520, 0.2068590, 0.1116020, -0.0059451, -0.0894573, 0.0617414, 0.1435130, 0.0796905, 0.0125305, 0.1085390, 0.0247227, -0.0277629, -0.0024571, -0.0003229, 0.0012920, 0.0103546, -0.0106631, -0.0164188, -0.0568550, 0.0814357, 0.0269486, -0.1084900, -0.1312440, -0.0582799, -0.1737650, -0.1614230, -0.1084430, -0.1222190, 0.0547736, 0.0218422, 0.1035710, 0.0505919, 0.0172878, 0.1239620, 0.0842178, 0.0065643, 0.1280380, 0.1073900, 0.0033204, -0.0505904, -0.0089756, -0.0004512, 0.0007733, 0.0088420, 0.0046793, -0.0745362, 0.0867803, -0.0288933, -0.0898602, -0.1502590, -0.0455147, -0.0503216, -0.0765177, -0.1034450, 0.0344278, 0.0892354, 0.0600338, 0.1526920, 0.1840780, -0.0668432, 0.2106850, 0.0314651, 0.0917470, 0.1516250, 0.1599450, 0.0597286, -0.0562202, -0.0456400, -0.0007958, -0.0009939, -0.0001021, -0.0059756, 0.0059784, -0.1118230, -0.1156010, -0.0295223, -0.0486842, -0.0676776, -0.0418525, -0.0477763, -0.1402360, -0.0615344, 0.1774690, 0.0716666, 0.0875325, -0.0136577, 0.0199230, -0.1230670, -0.0388063, -0.0305183, 0.0591164, 0.1687850, 0.0557864, -0.0905482, -0.0750084, -0.0004287, -0.0021150, 0.0001570, -0.0004730, -0.0298011, -0.0402610, -0.1746850, -0.1948710, -0.0762271, -0.1859970, 0.0100104, 0.0141201, -0.0622938, -0.0950794, 0.1562120, 0.0405879, 0.1078830, 0.1261290, 0.1046360, -0.0174896, 0.0889589, 0.0474537, -0.0515373, 0.0813138, -0.0744943, -0.0717250, -0.0936186, -0.0444926, -0.0427723, -0.0035386, -0.0002195, 0.0006087, -0.0325336, -0.0951248, -0.1684800, -0.1524870, -0.0364741, -0.1845130, -0.0957929, 0.0254724, 0.0736886, 0.1413140, 0.0382526, -0.1458960, 0.1215090, 0.0214734, 0.1577360, 0.0706191, 0.1519460, -0.0324796, -0.2222560, -0.0485154, 0.0112820, 0.0962036, 0.0518066, 0.0549371, -0.0092330, -0.0106889, -0.0007506, -0.0004864, -0.0048412, -0.0878337, -0.2129410, -0.2382620, -0.2094190, 0.0235527, 0.0458034, 0.0668059, -0.0421649, 0.1480100, -0.0571565, -0.0349147, 0.0603500, 0.1080350, -0.0681785, 0.1111850, -0.0295117, -0.1629920, -0.2659610, -0.0957737, 0.0463551, 0.1180560, 0.0327841, 0.0305466, -0.0030399, -0.0026610, 0.0002386, -0.0002915, -0.0020334, -0.0273103, -0.2076640, -0.2611830, -0.1460090, -0.0140140, -0.0036005, -0.0221827, 0.0293505, 0.0965633, -0.1817490, -0.0730674, 0.0356824, 0.1392200, 0.0053140, -0.0389051, -0.2184490, -0.1581750, -0.0966867, -0.0971920, -0.0688112, 0.0289225, -0.0425716, -0.0111752, -0.0014794, -0.0002943, 0.0002747, -0.0002694, -0.0034933, -0.0403083, -0.1096950, -0.3176500, -0.0881138, 0.0417062, -0.0558304, -0.1053110, -0.1244970, -0.0864638, -0.0600173, -0.0991870, 0.0108096, 0.0973347, 0.1477070, 0.0050927, 0.0448658, -0.0700960, -0.0826448, -0.0806831, -0.0461665, 0.0122476, -0.0856628, -0.0543442, -0.0008070, -0.0004491, 0.0003790, 0.0001805, -0.0047105, -0.0223951, -0.0364490, 0.0540679, 0.1183840, 0.1417220, 0.2007610, -0.0518821, -0.0669496, -0.0036837, -0.0570206, 0.0368226, -0.0216283, -0.0309799, 0.0519017, 0.0853929, -0.0738333, -0.1757540, 0.0094682, -0.0165018, -0.0800523, 0.0231095, 0.0036233, -0.0263544, 0.0006321, 0.0006996, -0.0002790, 0.0006154, 0.0005682, -0.0258020, 0.0293326, 0.1470070, 0.1084000, -0.0077538, 0.1534960, 0.1394860, -0.0098732, -0.0139355, -0.1278760, 0.0582982, -0.1863740, -0.0114817, 0.0433498, -0.0455971, -0.1169080, -0.0058821, -0.0736090, -0.0709483, -0.0807464, -0.1099060, -0.0353974, -0.0025672, 0.0083444, -0.0002610, -0.0000219, 0.0004906, -0.0063589, -0.0435964, -0.0490502, -0.0356928, -0.0509430, 0.0111657, 0.0109166, 0.0396625, 0.1332030, -0.0957493, -0.0085857, 0.0457823, -0.1557700, -0.1246830, -0.0348519, -0.0693903, -0.0997581, -0.0158861, -0.1263150, -0.1260530, -0.1406870, -0.1419620, -0.0784485, 0.0178957, 0.0088947, 0.0005972, 0.0000757, -0.0000196, -0.0079887, -0.0129567, -0.0468040, -0.0374206, -0.1315180, -0.1116230, -0.0516431, -0.0143117, -0.0163546, 0.0047835, 0.0603702, 0.3281290, 0.1504540, 0.0503262, 0.0671761, 0.0084153, 0.0184817, -0.1537120, -0.2056200, -0.1279210, -0.1163730, -0.0822051, -0.0366765, -0.0015442, 0.0000140, 0.0002774, 0.0002554, -0.0000816, -0.0019452, 0.0030543, -0.0265426, -0.0331130, -0.0933214, -0.0953786, 0.0157823, -0.0912639, -0.0913371, 0.0716800, 0.0861137, 0.0629052, 0.0565487, -0.0249400, 0.0419544, -0.0404942, -0.0745949, -0.2468560, -0.1708230, -0.1106010, -0.0481797, 0.0135830, -0.0036545, 0.0000869, 0.0005060, 0.0001490, 0.0001019, -0.0003215, 0.0004246, -0.0002209, -0.0016589, -0.0462476, -0.0743337, -0.0679151, -0.0720385, -0.0810903, -0.1314830, -0.1473480, -0.1723090, -0.1391910, -0.1182880, 0.0058996, 0.0481091, -0.0290945, -0.0273430, -0.0258332, -0.0547328, -0.0708932, -0.0268237, -0.0098079, -0.0017526, 0.0001125, 0.0002152, -0.0003248, -0.0002191, -0.0003299, -0.0001119, 0.0002347, 0.0005113, 0.0012863, 0.0000768, -0.0104565, -0.0076258, 0.0067648, 0.0143351, 0.0033226, 0.0089187, 0.0286165, -0.0142253, -0.0110749, -0.0029500, -0.0035345, -0.0403840, -0.0145956, -0.0054587, -0.0053104, -0.0132141, -0.0001621, -0.0002462, -0.0000518, 0.0003005, 0.0005547, 0.0005017, 0.0003417, 0.0005156, -0.0005799, -0.0003289, 0.0003080, 0.0002153, -0.0002026, -0.0005443, -0.0000155, -0.0002491, -0.0000362, 0.0008848, 0.0004049, -0.0002092, -0.0000238, -0.0001995, -0.0004874, -0.0003552, -0.0003460, 0.0000113, 0.0005768, -0.0005318, -0.0000948, -0.0003511, 0.0000383, 0.0001099, 0.0000532, -0.0004529, -0.0001624, 0.0004796, 0.0000320, 0.0001740, 0.0000467, 0.0003068, 0.0000069, -0.0000238, -0.0001619, -0.0016537, -0.0063152, -0.0002852, 0.0011523, 0.0087804, 0.0448993, 0.0334157, 0.0160667, 0.0046870, 0.0117603, 0.0187377, 0.0156275, 0.0012687, 0.0000278, 0.0002506, 0.0001123, -0.0000300, 0.0002314, -0.0000043, -0.0000965, -0.0000811, 0.0009823, 0.0014335, 0.0001440, 0.0002692, 0.0001640, -0.0005229, -0.0031788, -0.0215140, -0.0332750, 0.0096054, -0.0249847, -0.0396970, 0.0039847, 0.0026207, -0.0073925, 0.0748362, 0.0489993, 0.0174990, -0.0011929, -0.0007676, 0.0036706, 0.0017560, 0.0004104, 0.0001484, -0.0003306, -0.0003661, 0.0007411, 0.0002006, 0.0038785, 0.0037628, -0.0005562, -0.0012528, -0.0011835, -0.0231292, -0.0287376, -0.0309792, -0.1068680, -0.0504197, -0.0782426, -0.0509338, 0.0130941, -0.0150066, 0.0585860, 0.1713180, 0.0602553, 0.0579530, -0.0215167, 0.0056434, 0.0048402, -0.0022889, 0.0272559, 0.0081389, -0.0002473, -0.0003850, 0.0007205, 0.0000037, 0.0001276, 0.0031170, 0.0036788, -0.0030590, -0.0311929, -0.0992892, -0.2277340, -0.2860040, -0.2107680, -0.2315490, -0.1363720, -0.0187810, 0.0379730, 0.0573720, -0.0760982, -0.0856629, 0.0588856, -0.0055431, 0.0219984, 0.0934437, 0.1132700, 0.0694466, 0.0408566, 0.0122362, 0.0012939, 0.0001742, 0.0001716, -0.0002143, 0.0028698, 0.0545935, 0.1133830, 0.0686728, 0.0085953, -0.0619862, -0.0381337, -0.0898982, -0.1776430, -0.2120530, 0.1015030, 0.0716205, -0.0427944, -0.1482060, -0.0301596, -0.1442570, -0.0753183, 0.0576598, -0.1258830, -0.0494794, 0.0028584, 0.0442150, 0.0284218, 0.0164900, -0.0010766, 0.0005644, -0.0000432, 0.0012568, 0.0192511, 0.0769439, 0.0617554, 0.0281946, -0.0274883, -0.0700405, -0.1857980, -0.0524282, -0.2036400, -0.1536910, 0.0192214, -0.0518016, 0.0393519, 0.0554600, 0.0929111, 0.1703130, 0.1057390, 0.2013160, 0.0187339, -0.0493770, -0.0733107, -0.0047502, 0.0350211, 0.0256373, -0.0006927, 0.0000951, -0.0008204, -0.0033538, 0.0392777, 0.0419978, -0.0259616, -0.0637981, -0.0867003, -0.2724920, -0.2444630, -0.1365910, -0.2290580, 0.1503310, -0.1908370, -0.0905033, 0.0854404, 0.2828320, 0.3552940, 0.1678900, 0.1827300, 0.1946530, 0.0358451, 0.0039315, 0.0719386, -0.0745950, 0.0011671, 0.0274306, 0.0015518, 0.0015090, -0.0015635, 0.0053774, 0.0444339, 0.0022789, 0.0080412, -0.0233302, -0.0839905, -0.1994180, -0.2102080, -0.2116520, -0.2379260, -0.0850184, -0.1333760, -0.1326680, 0.1183300, 0.4423790, 0.3640090, 0.1984620, -0.0199276, 0.0297248, 0.1205210, 0.1107310, -0.0267557, 0.0074573, -0.0006575, 0.0416149, 0.0058837, 0.0003265, 0.0033472, 0.0059062, 0.0154411, 0.0337434, 0.0340231, 0.0185949, -0.1432860, -0.1053910, -0.1030680, -0.1395610, -0.1085750, 0.1165330, -0.0685289, -0.1559360, -0.0083870, 0.1482710, 0.2338760, 0.0065076, 0.0882311, 0.1040850, 0.0750237, 0.2003660, 0.0309338, 0.1164320, 0.1541700, 0.0460717, 0.0180476, 0.0004022, 0.0007973, 0.0215506, -0.0070523, 0.0717181, -0.0115780, -0.1115840, -0.1469990, -0.0883728, -0.1438380, -0.0145118, 0.1117780, -0.0372669, -0.0053898, 0.0186662, -0.0151516, 0.2069600, -0.0097955, 0.1197930, 0.1829240, 0.2469160, 0.0280067, 0.2262600, 0.1849240, 0.1631070, 0.0940779, 0.0083726, 0.0032828, 0.0003528, 0.0032978, 0.0165420, 0.0007371, 0.0124750, -0.0531904, -0.1010700, 0.0492094, -0.0462765, -0.1243920, -0.0025783, -0.0172913, -0.1748070, 0.1309550, 0.2766660, 0.0265647, -0.0764470, 0.1882590, 0.2928750, 0.2552080, 0.3012690, 0.2375540, 0.1964010, 0.1900410, 0.1676910, 0.0166030, 0.0125277, 0.0015314, -0.0000888, 0.0003142, 0.0043521, 0.0017417, -0.0153591, -0.0454617, -0.0972373, -0.0916195, -0.1882540, 0.0140081, -0.0175148, -0.0716265, -0.2756710, -0.1465130, 0.2734660, 0.1532760, -0.1043600, 0.0179967, 0.1595770, 0.1491590, 0.0009187, -0.1258110, 0.0901275, 0.1842600, -0.0163937, -0.0266343, 0.0095632, 0.0036485, 0.0005293, -0.0001503, 0.0013842, 0.0046433, 0.0632242, -0.0517690, -0.1577180, -0.2196990, -0.1031490, -0.0569945, -0.1367410, -0.1422990, -0.1751280, -0.0653755, 0.1310640, 0.0833074, -0.0470368, -0.1310010, -0.1609580, -0.0904492, -0.1136490, -0.0919171, -0.0271961, -0.0774207, -0.0835079, -0.0350975, -0.0225090, -0.0030900, 0.0002240, 0.0010612, 0.0001466, 0.0064878, 0.0086235, -0.0368759, -0.0722270, -0.1748210, -0.0543359, -0.1652430, -0.0341593, -0.2289210, -0.2613350, -0.0576424, 0.0348660, 0.0440127, -0.2284620, -0.2461160, -0.2726630, -0.1127890, 0.0460345, -0.0307470, -0.2324520, -0.1705740, -0.0741004, -0.0577297, -0.0114036, -0.0001884, -0.0002182, 0.0004218, -0.0045453, -0.0505959, 0.0366973, 0.0346020, 0.1157000, 0.1075580, -0.1336870, -0.2767180, -0.0373944, -0.1780870, -0.1079740, -0.0752217, -0.0740654, 0.1312290, -0.0390551, -0.1316060, -0.1701290, -0.1037890, -0.1026570, -0.2761280, -0.2033650, -0.0871825, -0.0811728, -0.0581286, -0.0198657, -0.0039295, 0.0003116, 0.0007488, -0.0160391, -0.0824786, 0.0661951, 0.1217300, 0.1549450, -0.0269492, -0.0684621, -0.0918685, 0.0919643, -0.2209800, -0.1025780, -0.1168660, -0.2745330, -0.0911390, 0.1747660, -0.1485390, -0.1510300, -0.1332750, -0.2422400, -0.4066150, -0.2736420, -0.2472390, -0.0983226, -0.0653812, -0.0202670, -0.0019405, 0.0007615, 0.0000556, -0.0411603, -0.0790447, -0.0611755, 0.0371314, -0.0218837, 0.0741209, -0.0946739, -0.0266463, -0.0687393, -0.0676540, -0.0439938, -0.1281180, -0.0152750, 0.0401833, 0.3409900, 0.1735750, -0.0077868, -0.1368260, -0.3555340, -0.4474650, -0.2647700, -0.0837455, -0.0323890, -0.0093414, -0.0003000, 0.0034934, 0.0020195, 0.0001020, -0.0113652, -0.1255090, -0.0942642, 0.0438403, -0.1168460, -0.0631393, -0.0984136, -0.0157351, 0.0042044, 0.1948170, 0.0701502, 0.0271352, 0.0024219, 0.2316930, 0.4222540, 0.3713020, 0.0465020, -0.4545460, -0.5087490, -0.4268030, -0.2510450, -0.1740120, -0.0937996, 0.0003356, 0.0018239, -0.0031458, -0.0000154, 0.0130576, 0.0101637, -0.0705998, -0.1049480, 0.0056424, 0.0551895, -0.0408438, -0.0521595, -0.0393593, -0.0083495, -0.0510184, 0.1000240, 0.0028206, 0.1309820, 0.0648546, 0.2699960, 0.3166940, -0.0836456, -0.6341840, -0.4372990, -0.2974070, -0.1514620, -0.1006770, 0.0097033, 0.0319331, -0.0062322, -0.0007719, 0.0000388, 0.0047803, 0.0014365, -0.0493511, -0.1017720, -0.0378380, 0.0623866, -0.1078000, -0.0128991, 0.0145021, 0.1347020, 0.0556604, 0.0574085, 0.1091950, -0.0369700, 0.0784687, 0.0277079, 0.2193850, -0.5216880, -0.8209180, -0.5295420, -0.2371090, -0.0593632, -0.0714507, 0.0126953, 0.0151494, -0.0036670, -0.0000233, 0.0003118, -0.0005654, -0.0074893, -0.0514320, -0.1726690, -0.1969270, -0.0189953, 0.0328367, 0.0380959, 0.0156400, 0.0724502, -0.0442976, -0.0389969, -0.1818740, -0.0147908, 0.0000416, -0.1401650, -0.2048130, -0.6952940, -0.6081020, -0.3082100, -0.1093220, -0.0586622, -0.0377498, -0.0161735, -0.0003245, 0.0059131, 0.0003303, 0.0002252, 0.0000185, -0.0071507, -0.0424889, -0.1251670, -0.1659400, 0.0728233, 0.0217709, -0.0383419, 0.1296900, 0.0720792, -0.0002758, 0.0869950, 0.1339810, 0.1771920, -0.0641624, -0.2432310, -0.5090030, -0.6462850, -0.3856790, -0.1861360, -0.0872939, -0.0215227, -0.0079253, -0.0071762, -0.0077304, -0.0022748, 0.0001757, 0.0004636, 0.0002562, 0.0012354, -0.0093115, -0.0188440, -0.0078165, -0.0382975, 0.0053321, -0.1098470, -0.1335190, -0.0967593, 0.0395086, 0.0659783, -0.0610230, -0.1293260, -0.1762520, -0.5777800, -0.5844370, -0.4288580, -0.3041000, -0.1356410, -0.1054620, -0.0277775, -0.0367365, 0.0036672, -0.0076362, -0.0062262, -0.0000176, -0.0004581, 0.0001400, 0.0039448, 0.0197126, 0.0661912, 0.2323610, 0.1613970, 0.1392790, 0.1627480, -0.0189697, 0.1808900, 0.0530323, 0.2090690, 0.0932897, 0.0769679, -0.0810485, -0.4028830, -0.4501940, -0.4208640, -0.2622330, -0.1665930, -0.1894550, -0.1192270, -0.0306179, -0.0062552, -0.0079740, -0.0013137, -0.0002676, -0.0004113, -0.0001796, 0.0001443, 0.0027101, 0.0380178, 0.0923027, 0.0851851, 0.1195410, 0.2461860, 0.2833790, 0.0766458, 0.0325695, 0.1307470, 0.2063850, 0.0850007, -0.0858265, -0.1137530, -0.2135270, -0.2019170, -0.1082110, -0.0698638, -0.0322386, 0.0012942, -0.0065671, -0.0023939, -0.0008322, -0.0011299, -0.0003631, -0.0003712, -0.0003341, -0.0002613, 0.0003114, -0.0002601, 0.0091853, 0.0441857, 0.0785105, 0.0890266, 0.1390410, 0.1214110, 0.1789940, 0.1593280, 0.2249160, 0.2119950, 0.1189720, 0.0375600, 0.0017869, 0.0275453, 0.0170713, 0.0022804, 0.0039419, 0.0061785, -0.0010427, 0.0000318, -0.0000101, -0.0001521, 0.0005248, -0.0009239, 0.0003836, -0.0002144, -0.0002982, 0.0002934, -0.0006532, 0.0039455, 0.0191656, 0.0168321, 0.0024106, 0.0080776, 0.0057343, 0.0053138, -0.0039337, 0.0333090, 0.0096618, 0.0065617, 0.0095448, 0.0284432, 0.0018409, 0.0003654, 0.0012231, 0.0039646, 0.0003290, -0.0003470, -0.0002399, -0.0002014, 0.0001640, -0.0007066, 0.0001878, 0.0001781, -0.0001053, -0.0003886, -0.0002616, -0.0005062, -0.0005816, 0.0000362, 0.0002207, 0.0003250, 0.0004926, -0.0003421, -0.0007278, 0.0001700, -0.0004090, 0.0005564, -0.0000475, -0.0000435, -0.0004103, -0.0005314, -0.0003147, -0.0008800, 0.0004864, 0.0000641, 0.0000023, 0.0002309, -0.0007615, 0.0002099, -0.0005068, -0.0001642, -0.0005044, -0.0003498, -0.0004657, -0.0006023, -0.0013852, -0.0043297, -0.0034118, -0.0107479, -0.0103300, -0.0164846, -0.0261771, -0.0148594, -0.0125921, -0.0191536, -0.0138407, -0.0101593, -0.0154565, -0.0249597, -0.0096902, -0.0026899, -0.0008217, 0.0002758, 0.0002166, -0.0001142, 0.0001204, 0.0002283, 0.0001243, 0.0000401, 0.0003388, -0.0019356, -0.0007567, -0.0032674, -0.0081871, -0.0132180, 0.0093207, -0.0021292, -0.0488547, -0.0408094, -0.0238968, -0.0890838, -0.0766542, -0.1173970, -0.1639330, -0.1483850, -0.1094830, -0.0787463, -0.0567282, -0.0205074, -0.0044174, 0.0073355, 0.0061776, 0.0000724, -0.0005498, 0.0002082, 0.0001161, 0.0050265, -0.0000887, -0.0022995, 0.0243547, 0.0097781, 0.0169161, 0.0208623, -0.0549161, -0.0575274, 0.0465681, 0.1438070, 0.1108860, -0.1486920, -0.1414960, -0.1714670, -0.3341680, -0.3640020, -0.2723300, -0.1882810, -0.1328850, -0.0534103, -0.0164193, 0.0001228, 0.0012326, -0.0045641, -0.0003942, 0.0002099, -0.0004327, 0.0142619, 0.0041851, 0.0057807, 0.1159730, 0.1696950, 0.1200670, 0.2177880, 0.0478740, 0.1268400, 0.0775592, 0.1267580, 0.0625014, -0.0453947, 0.0106894, -0.1445510, -0.3154090, -0.2842740, -0.3796680, -0.3429860, -0.2329670, -0.1260100, -0.0895413, -0.0596229, -0.0211336, -0.0026709, 0.0003162, 0.0004185, 0.0001815, 0.0026642, 0.0202133, 0.0938610, 0.2080350, 0.2278590, 0.1970210, 0.1471060, 0.0927077, -0.0836438, 0.0308996, 0.2900310, 0.1189230, 0.0487551, 0.1594970, 0.0325350, -0.0951297, -0.2171900, -0.5155130, -0.6563120, -0.4234280, -0.1991480, -0.1591460, -0.0619745, -0.0183972, -0.0049914, -0.0016176, 0.0000100, -0.0001699, 0.0021232, 0.0769029, 0.1797470, 0.1454550, 0.2269510, 0.1156070, -0.1038250, 0.0598274, 0.0202623, 0.0675251, -0.0188549, 0.1762570, 0.0764613, -0.0425260, 0.0978502, -0.0742053, -0.0171886, -0.3676770, -0.3737700, -0.3661760, -0.3023720, -0.1575550, -0.0686033, -0.0354096, -0.0147910, -0.0054960, -0.0003485, 0.0050998, 0.0005606, 0.1387010, 0.2618060, 0.0564988, 0.1077740, 0.0434373, -0.1040940, -0.0634260, 0.0151093, -0.0206121, -0.1561010, 0.1233920, 0.0490104, 0.1167740, 0.0263441, -0.1123130, -0.1265820, -0.2071110, -0.4399230, -0.5579820, -0.4242900, -0.2397920, -0.1552060, -0.0354514, -0.0091113, -0.0009117, -0.0003721, 0.0014476, 0.0039622, 0.0438888, 0.2508390, 0.0082545, -0.0828309, -0.1082400, -0.2777830, -0.1117400, 0.3038790, -0.2140120, 0.0681528, 0.2399080, 0.1324390, 0.1451940, 0.1813910, 0.1212890, -0.0250379, -0.1944800, -0.6497980, -0.6414770, -0.3904490, -0.2367780, -0.1703610, -0.0482952, -0.0020202, -0.0037291, 0.0000250, 0.0021696, 0.0052166, 0.0330731, 0.1593100, 0.1458190, -0.0031047, -0.1192940, -0.2772970, -0.1101070, -0.2028640, -0.1596710, 0.2854570, 0.2407510, 0.3696650, 0.5816680, 0.6006470, 0.1969810, -0.2672140, -0.4279400, -0.7105010, -0.5364120, -0.2862940, -0.1200300, -0.0537666, -0.0223378, -0.0050641, 0.0072600, 0.0000602, 0.0019560, 0.0063499, 0.0355754, 0.0537454, 0.1084130, 0.0137019, -0.1706000, -0.4330400, -0.3066030, -0.0481525, 0.0531931, -0.0062665, 0.2241220, 0.4519930, 0.5315640, 0.5945810, 0.1478620, -0.3050620, -0.4375080, -0.4895800, -0.3959160, -0.0941555, -0.0046896, -0.0828901, -0.0548064, -0.0028353, 0.0071373, 0.0002295, 0.0041363, 0.0128936, 0.0671394, 0.0655586, -0.0203770, -0.0499043, -0.1985530, -0.0454129, 0.0125162, -0.0180857, 0.3283770, 0.2865200, 0.3544880, 0.4444490, 0.3562590, 0.0408356, -0.4804030, -0.6821840, -0.5035640, -0.3109240, -0.2394140, 0.0479768, 0.1080470, -0.0302356, -0.0435688, -0.0071697, 0.0021626, -0.0002162, 0.0027640, 0.0075768, 0.0030059, -0.0229441, -0.0001393, -0.2001730, -0.2023790, -0.1424840, 0.0139318, 0.0813351, 0.0226751, 0.0438079, 0.0834424, 0.3932460, 0.2452920, -0.0197894, -0.3721670, -0.2797350, -0.2225900, -0.1343140, 0.0312103, 0.1825740, 0.1669360, 0.1345510, 0.1049960, -0.0060047, 0.0099861, 0.0008652, 0.0008288, 0.0024115, -0.0179065, -0.0688598, -0.1150300, -0.1341950, -0.1432630, -0.2070340, -0.1170400, -0.0615721, 0.1199440, 0.0141827, 0.1215990, 0.2562730, 0.1800720, 0.1156560, -0.1519250, 0.0450205, -0.0110277, 0.0734471, 0.0860318, 0.0970314, 0.0889713, 0.1528310, 0.1481980, 0.0573946, 0.0172386, -0.0008912, -0.0000021, 0.0003821, -0.0118698, -0.0623290, -0.0685107, -0.1038750, -0.2041460, -0.1071280, -0.1346340, -0.0675979, -0.0665138, -0.1162950, 0.0142157, 0.1022410, 0.1298410, -0.1323390, -0.2727790, -0.1551050, 0.1266250, 0.0929832, 0.2292540, 0.0688824, 0.0454903, -0.0117393, 0.1228660, 0.0546403, 0.0010215, -0.0003924, -0.0004034, 0.0003221, 0.0338098, -0.0874360, -0.0757154, 0.0270597, 0.0858976, 0.2303320, -0.0181092, -0.0632188, -0.0277747, -0.1428640, 0.1797530, 0.1672290, 0.2272780, -0.0407641, -0.0071199, -0.1403850, 0.0657331, 0.2053140, 0.1258630, 0.2758300, 0.1012100, 0.0833045, 0.0576493, 0.0897147, 0.0115630, 0.0003604, 0.0004986, -0.0004543, 0.0260027, -0.0617183, -0.1136530, 0.0541767, 0.3259960, 0.1953430, 0.2918990, -0.0155198, -0.1435190, -0.1061180, -0.0170525, 0.2526370, -0.0268704, -0.2008290, -0.2117790, 0.0714046, -0.0187616, -0.0013667, 0.0253697, 0.1350000, 0.1422060, 0.1768780, 0.0402485, 0.1244040, 0.0242898, -0.0000558, -0.0000472, 0.0006448, -0.0154115, -0.0711613, -0.1725450, 0.0195381, 0.1106220, -0.0873376, -0.0227855, -0.1684040, -0.2160890, -0.1557340, -0.0283050, 0.1239570, -0.1590810, -0.1127290, -0.0163808, -0.0139170, 0.0508679, -0.0101584, 0.1488100, 0.1564930, 0.1128630, 0.1665500, 0.0857429, 0.0462664, 0.0061601, 0.0016705, 0.0003365, -0.0002011, -0.0179314, -0.0220794, -0.0941638, -0.0655182, -0.1993970, -0.1027800, -0.0312848, 0.0977680, 0.0117110, -0.1496190, -0.0669796, -0.2234640, -0.1545460, -0.0623073, 0.0589438, 0.0285173, 0.1561030, 0.1319780, 0.1229940, 0.2698920, 0.1940330, 0.1534000, 0.0794330, 0.0105782, 0.0058137, 0.0000995, -0.0022271, -0.0581662, -0.0703254, -0.0069122, -0.0515867, -0.3143860, -0.1659190, -0.1319790, -0.0510441, 0.0029781, -0.1886610, -0.1806860, -0.0301084, 0.0460746, -0.1134940, 0.0554554, 0.0540202, 0.0821923, 0.1341280, 0.1999690, 0.0162622, 0.1443060, 0.0940426, 0.0250580, 0.0473722, 0.0281785, 0.0016112, 0.0002284, -0.0053676, -0.0496818, -0.0628296, -0.0861603, -0.1258000, -0.0736600, 0.0766817, 0.0616148, 0.1343790, -0.0500499, -0.1097640, -0.1247700, -0.0643484, 0.0007026, -0.2889970, -0.0716935, -0.1275010, 0.0125131, -0.0673526, 0.0588380, -0.0345651, -0.0527153, 0.0281442, -0.0569541, -0.0630114, 0.0079139, -0.0003358, 0.0000671, 0.0003586, 0.0052504, 0.0029209, -0.0910388, -0.1887040, -0.1519330, -0.1502980, -0.1044120, -0.0676384, -0.0908218, -0.0547860, -0.1012660, -0.2866530, -0.0755560, -0.0474645, 0.0304731, -0.1347440, -0.0761485, -0.0288124, -0.1766800, -0.1723190, -0.0607643, -0.0557320, -0.1358480, -0.0718046, -0.0002833, -0.0000091, -0.0003117, -0.0003556, 0.0034803, 0.0172027, 0.0155366, -0.1048760, 0.0035633, -0.1029860, -0.1571740, -0.1552900, -0.0153199, -0.1870220, -0.1527220, -0.0541923, -0.1970850, -0.1225000, -0.2421660, -0.1914780, 0.0674154, 0.0339835, 0.0663204, 0.0421276, 0.0018587, -0.1486480, -0.1382050, -0.0699673, -0.0086210, 0.0002301, 0.0001539, 0.0002668, 0.0031386, 0.0157671, 0.0271898, -0.0338912, -0.0853320, -0.0171999, -0.0667554, 0.0357815, -0.0013014, 0.0732599, -0.1249300, 0.0901337, -0.2486330, -0.0562081, -0.2112980, 0.0233428, -0.0440982, -0.1513900, 0.0655051, -0.0000644, -0.0635499, -0.1544310, -0.1218790, -0.0460691, -0.0045075, -0.0003013))
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s1,
    done => done_s2,
    start => start_s3,
    ack => ack_s4,
    in_a => in_a_s5,
    out_a => out_a_s6,
    out_offset => out_offset_s7,
    op_argument => op_argument_s8,
    op_result => op_result_s9,
    op_send => op_send_s10,
    op_receive => op_receive_s11
);
interlayer_u13 : interlayer generic map(
    width => 56,
    word_size => 9
) port map(
    clk => clk,
    rst => rst,
    ready => ready_s14,
    done => done_s15,
    start => start_s16,
    ack => ack_s17,
    previous_a => previous_a_s18,
    next_a => next_a_s19
);

in_a_s5 <= next_a_s19;
start_s3 <= start_s16;
ready_s14 <= ready_s1;
op_result_s9 <= resize(op_argument_s8, mk(fixed_spec(fixed_spec'(int => 2, frac => 8))));

uPS : ps port map(
    clk => clk,
    rst => rst_sink
);
previous_a_s18 <= to_vec(reals'(0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.3176470, 0.9882350, 0.9882350, 0.9882350, 0.9882350, 0.9882350, 0.9882350, 0.9921570, 0.9882350, 0.9882350, 0.9882350, 0.7254900, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.1411760, 0.6196080, 0.9176470, 0.5725490, 0.7176470, 0.7725490, 0.7490200, 0.9921570, 0.9921570, 0.9921570, 0.9921570, 0.5058820, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000, 0.0000000));
done_s15 <= start;
test_out <= shift_range(std_logic_vector(get(out_a_s6, to_integer(sel), mk(fixed_spec(fixed_spec'(int => 2, frac => 8))))), 8)(test_out'range) when to_integer(sel) < 40 else "00000000";
end system;
