library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package fc_weights_defs is
end fc_weights_defs;

package body fc_weights_defs is
end fc_weights_defs;